// load_tableをノンブロッキング代入すべきかは要調査。

`default_nettype none
module sqrt_load_const_table (
    input wire [9:0] addr,
    output wire [81:0] cst,
    input wire clk,
	input wire rstn);

(* RAM_STYLE="BLOCK" *) reg [81:0] ram [1023:0];
//always @(posedge clk)
//    cst <= ram[addr];
assign cst = ram[addr];
initial begin
	ram[0] = 82'b1011010100000100111100100010010011011101001001111110111011000001101000110000000000;
	ram[1] = 82'b1011010011101110010101011100010001100010011000100100111010001111010001001001101011;
	ram[2] = 82'b1011010011010111110000011101101011000001101110111110001110110100111100100100110110;
	ram[3] = 82'b1011010011000001001101100110001011100101010111010111100100110001111101001110111000;
	ram[4] = 82'b1011010010101010101100110101011101011100010011000010111100101111101101010101100100;
	ram[5] = 82'b1011010010010100001110001011001100011001110000101111010010010000001111010011111011;
	ram[6] = 82'b1011010001111101110001100111000010110101111111110101110000100010100101111000111110;
	ram[7] = 82'b1011010001100111010111001000101011111101100110001101111001011100000000010001001101;
	ram[8] = 82'b1011010001010000111110101111110011000001101010001010101011111010000001000010001000;
	ram[9] = 82'b1011010000111010101000011100000100000111010100110000111110100111111000110110011000;
	ram[10] = 82'b1011010000100100010100001101001010101000100001011101001100100101010000110111010000;
	ram[11] = 82'b1011010000001110000010000010110000100100101111101100000000110010101001001111001101;
	ram[12] = 82'b1011001111110111110001111100100010111101111001000000100110011101010110101010000100;
	ram[13] = 82'b1011001111100001100011111010001100101011110101110111100000010111110111011111101011;
	ram[14] = 82'b1011001111001011010111111011011001011010010111101001001111001001111010010101011010;
	ram[15] = 82'b1011001110110101001101111111110100111001100111101111010100011011110101001110101001;
	ram[16] = 82'b1011001110011111000110000111001011101101010100111000111110100101010111010010000000;
	ram[17] = 82'b1011001110001001000000010001001000001111110101111000000100110111111100011001011000;
	ram[18] = 82'b1011001101110010111100011101010111111100101111001100000100001010000010110101110010;
	ram[19] = 82'b1011001101011100111010101011100110000110010000100000101011000110000011000111000000;
	ram[20] = 82'b1011001101000110111010111011011110110010001010001000000111110101011011001110101100;
	ram[21] = 82'b1011001100110000111101001100101110001010011101010001011111001111101011100010101000;
	ram[22] = 82'b1011001100011011000001011111000001001100010111111001001001101011100101000010000000;
	ram[23] = 82'b1011001100000101000111110010000010101100011101001011011000110010000100111111111001;
	ram[24] = 82'b1011001011101111010000000101011111110000011001111000001101101010000011000111000000;
	ram[25] = 82'b1011001011011001011010011001000100110011000111011110010000010000001101010111011101;
	ram[26] = 82'b1011001011000011100110101100011110010011101010101000011000110111001001010000000000;
	ram[27] = 82'b1011001010101101110100111111011001100100000000101011101000110011001001110101111000;
	ram[28] = 82'b1011001010011000000101010001100001101110000001010010000010111001001001000010101100;
	ram[29] = 82'b1011001010000010010111100010100100001011111101000101010001000000101010011000000000;
	ram[30] = 82'b1011001001101100101011110010001101101101011010000100000110100000000111100001101010;
	ram[31] = 82'b1011001001010111000010000000001010010111100000100100110110000010011110011001001001;
	ram[32] = 82'b1011001001000001011010001100001000011111001001110101101010111010110011000100000000;
	ram[33] = 82'b1011001000101011110100010101110100010001100010110000011100000011110101110101101101;
	ram[34] = 82'b1011001000010110010000011100111010000000000110010001111110011101101110111100100010;
	ram[35] = 82'b1011001000000000101110100001000111011101001011000010000000000000101000111100010111;
	ram[36] = 82'b1011000111101011001110100010001001110000100111100101110111100010100100111000100100;
	ram[37] = 82'b1011000111010101110000011111101110000110010001010101010000000010000001011010100001;
	ram[38] = 82'b1011000111000000010100011001100000111111101011111011001110101101011010110000110000;
	ram[39] = 82'b1011000110101010111010001111010000011110111100011110011010011000000000011100000001;
	ram[40] = 82'b1011000110010101100010000000101001111011101110111000000111001110101111101000000000;
	ram[41] = 82'b1011000110000000001011101101011010110001101001011010011100100000011110000010010001;
	ram[42] = 82'b1011000101101010110111010101001111110010000111001111011000010100100110110011000110;
	ram[43] = 82'b1011000101010101100100110111110111001110101011000110100000110110001100001000000111;
	ram[44] = 82'b1011000101000000010100010100111110101110100100111001010010110100011111000111000100;
	ram[45] = 82'b1011000100101011000101101100010011001110111110100001100100101010110001001101101000;
	ram[46] = 82'b1011000100010101111000111101100011001100110101101011010111111010110000010100001110;
	ram[47] = 82'b1011000100000000101110001000011100011010111010010011011011111101101001101000000000;
	ram[48] = 82'b1011000011101011100101001100101100000001111100000000001000110100111010000000000000;
	ram[49] = 82'b1011000011010110011110001001111111111100011000101010111101001000101100110001100001;
	ram[50] = 82'b1011000011000001011001000000000110110110001110000101001011001011100011010010010000;
	ram[51] = 82'b1011000010101100010101101110101110110001010011110100111111100011110110100101001001;
	ram[52] = 82'b1011000010010111010100010101100101000101100111001011000111010000000101010111000100;
	ram[53] = 82'b1011000010000010010100110100011000101010001011110110101011010011001100110011100011;
	ram[54] = 82'b1011000001101101010111001010110110111110100000010011110000001101101100001101110000;
	ram[55] = 82'b1011000001011000011011011000101111000000111100001110001010011001010011100011011011;
	ram[56] = 82'b1011000001000011100001011101101110011000011011010011100101011001111001011001111000;
	ram[57] = 82'b1011000000101110101001011001100011011101001001110111010000100011111111110100011000;
	ram[58] = 82'b1011000000011001110011001011111101011000010110011100100100001100010101011001101110;
	ram[59] = 82'b1011000000000100111110110100101001111100000000110100100100110110001101010101100011;
	ram[60] = 82'b1010111111110000001100010011011000011000100010001000001000100111001001000110000100;
	ram[61] = 82'b1010111111011011011011100111110110100111001101010110101100000101110001011001011000;
	ram[62] = 82'b1010111111000110101100110001110011010010010100000010011101000011100101010101010000;
	ram[63] = 82'b1010111110110001111111110000111101110100110111101001010100011100101011000101101000;
	ram[64] = 82'b1010111110011101010100100101000011100101111000000101000000000000000000000000000000;
	ram[65] = 82'b1010111110001000101011001101110101100001101100101010100001111000111010110100100001;
	ram[66] = 82'b1010111101110100000011101011000000011001011000011000101000101000001100011110000000;
	ram[67] = 82'b1010111101011111011101111100010100100011000100000101111110111101101101100000001101;
	ram[68] = 82'b1010111101001010111010000001100000010001001000010001001001100011101000011101001100;
	ram[69] = 82'b1010111100110110010111111010010010100110100010101010111101100011011000000000000000;
	ram[70] = 82'b1010111100100001110111100110011010101001101110111101000111111010100100100011010000;
	ram[71] = 82'b1010111100001101011001000101101000010001011100101001000100101001000100011011000000;
	ram[72] = 82'b1010111011111000111100010111101001111110000100111001010100111101101111000110011000;
	ram[73] = 82'b1010111011100100100001011100001110010011100111001010010111111111011110101011000000;
	ram[74] = 82'b1010111011010000001000010011000101111111110011010001000101100101101111101100010010;
	ram[75] = 82'b1010111010111011110000111011111111101101011001101100010010101110100001000011011101;
	ram[76] = 82'b1010111010100111011011010110101011100100000001000110111110111011110000000100101100;
	ram[77] = 82'b1010111010010011000111100010110111101000101000100111001001101001001001001010011001;
	ram[78] = 82'b1010111001111110110101100000010100001001100111110011111100011000010110001010110000;
	ram[79] = 82'b1010111001101010100101001110110001011000100010010010111100111011101111011101011001;
	ram[80] = 82'b1010111001010110010110101101111101100100101000101010110111111101111110110110000000;
	ram[81] = 82'b1010111001000010001001111101101001110010100110110110100010011111001111000111000101;
	ram[82] = 82'b1010111000101101111110111101100100011000011111100110010110011111000101001010110000;
	ram[83] = 82'b1010111000011001110101101101011110100001011010010110110111101101111100000111100101;
	ram[84] = 82'b1010111000000101101110001101000110101010001000011100010100111101011001010110100000;
	ram[85] = 82'b1010110111110001101000011100001110000100001001011011111101000101000110100000100001;
	ram[86] = 82'b1010110111011101100100011010100011010010111001111010100011001110001010101000110000;
	ram[87] = 82'b1010110111001001100010000111110111000010000001000001011111001111011111001000000000;
	ram[88] = 82'b1010110110110101100001100011111001010011111111101110100111011110100000010101101000;
	ram[89] = 82'b1010110110100001100010101110011010111010101100101000000010101111000100101001111000;
	ram[90] = 82'b1010110110001101100101100111001010100110101111110111110011111001101011000011100110;
	ram[91] = 82'b1010110101111001101010001101111000100100010111111100011011010000101000110001111000;
	ram[92] = 82'b1010110101100101110000100010010110011010111111010000101010110001010001000000001100;
	ram[93] = 82'b1010110101010001111000100100010011110000111100000010100001100111010111010011010101;
	ram[94] = 82'b1010110100111110000010010011100000001111111000011101011101110011011010100001100010;
	ram[95] = 82'b1010110100101010001101101111101100111100100010101100000010110111110001111011001000;
	ram[96] = 82'b1010110100010110011010111000101010010010110000011110000001100010001010100100000000;
	ram[97] = 82'b1010110100000010101001101110001000110001011110010110101000110101011110000110000111;
	ram[98] = 82'b1010110011101110111010001111111000001110111101101000001111011100101000110110010000;
	ram[99] = 82'b1010110011011011001100011101101001111100001100110001101001001011011001111000001000;
	ram[100] = 82'b1010110011000111100000010111001110100001011000101001011000011011111011111001001100;
	ram[101] = 82'b1010110010110011110101111100010110101001110001101000110010101001101100011010101101;
	ram[102] = 82'b1010110010100000001101001100110010011000000011010100001101000000001110000010010110;
	ram[103] = 82'b1010110010001100100110001000010011110100110101010010101001011100110110110001010111;
	ram[104] = 82'b1010110001111001000000101110101001110001101111010100101000101101011011101000000000;
	ram[105] = 82'b1010110001100101011100111111100111001000111000010000011110010001001111011100000111;
	ram[106] = 82'b1010110001010001111010111010111011011101100101001000111111011001000011100010000000;
	ram[107] = 82'b1010110000111110011010100000010111101101010100000111110001010000000011110000011001;
	ram[108] = 82'b1010110000101010111011101111101110001111010011010000110011110110111001000111100000;
	ram[109] = 82'b1010110000010111011110101000101110000100101011001000011010111011000010000011000000;
	ram[110] = 82'b1010110000000100000011001011001010010101110101110011110111001000100011010111010000;
	ram[111] = 82'b1010101111110000101001010110110010110101010100101101001101011001110100010110011000;
	ram[112] = 82'b1010101111011101010001001011011000101111010110010101010000000110100110000000000000;
	ram[113] = 82'b1010101111001001111010101000101110101001011101001001100111100001110010100101111000;
	ram[114] = 82'b1010101110110110100101101110100011110011111111001101110011011001010011110011101110;
	ram[115] = 82'b1010101110100011010010011100101010111010001111001010110100101110000100011101001011;
	ram[116] = 82'b1010101110010000000000110010110101010011111010100100000011000100100111101100000000;
	ram[117] = 82'b1010101101111100110000110000110011110000100011011100110001111111000110000001011101;
	ram[118] = 82'b1010101101101001100010010110011000011000101101100001110111010110000000111110101010;
	ram[119] = 82'b1010101101010110010101100011010100000001101101001110101101101111100010001111001001;
	ram[120] = 82'b1010101101000011001010010111011000001110110001100100110111110001010000000010111000;
	ram[121] = 82'b1010101100110000000000110010010111010000110111100110011001010000011111100011000000;
	ram[122] = 82'b1010101100011100111000110100000010000101111001001111101111011100000100000000101010;
	ram[123] = 82'b1010101100001001110010011100001011000100010110100100000101001111101000111101000101;
	ram[124] = 82'b1010101011110110101101101010100011001111110100001111110101111110010011110111000100;
	ram[125] = 82'b1010101011100011101010011110111101000100010010000101000010111001000110111000000000;
	ram[126] = 82'b1010101011010000101000111001001001000000001111111011111101000110011110110010000000;
	ram[127] = 82'b1010101010111101101000111000111010111010100111100110111100010010101111101000000000;
	ram[128] = 82'b1010101010101010101010011110000010101100110011010111001010010111100111001110000000;
	ram[129] = 82'b1010101010010111101101101000010011101000010111100110001110011000101100000010111111;
	ram[130] = 82'b1010101010000100110010010111011111000001101001010100110000001111100010010111110010;
	ram[131] = 82'b1010101001110001111000101011010110111010010110000101100111110001000101011110111111;
	ram[132] = 82'b1010101001011111000000100011101110000001010111111111000000000111010110010110100000;
	ram[133] = 82'b1010101001001100001010000000010101110011010010011010000101101011100110101101000101;
	ram[134] = 82'b1010101000111001010101000001000000011001111000101001101111001100011000110010110000;
	ram[135] = 82'b1010101000100110100001100101100000000001101000111111101100001010110001100100100011;
	ram[136] = 82'b1010101000010011101111101101100111100100000010011010000100110101000101101110001000;
	ram[137] = 82'b1010101000000000111111011001001000101000011100111101101011010100011010000110010111;
	ram[138] = 82'b1010100111101110010000100111110101100011010100110010101100010011000000010011000110;
	ram[139] = 82'b1010100111011011100011011001100000101011101110011100000111010111111101000110010011;
	ram[140] = 82'b1010100111001000110111101101111100011011010110001111110101000101111001111000011100;
	ram[141] = 82'b1010100110110110001101100100111011111000101010010100000110111111000010010010001000;
	ram[142] = 82'b1010100110100011100100111110010000111000010101110101001111101110110001111100111110;
	ram[143] = 82'b1010100110010000111101111001101101010001110011111011100001111010101010100010100101;
	ram[144] = 82'b1010100101111110011000010111000100111101010111010110010010010110110000000110000000;
	ram[145] = 82'b1010100101101011110100010110001001110111100010100011011000110110100000010000011011;
	ram[146] = 82'b1010100101011001010001110110101110101001100011111001101000011001001010010011010000;
	ram[147] = 82'b1010100101000110110000111000100101111111001101001001011100101001001110111010111001;
	ram[148] = 82'b1010100100110100010001011011100011010000101101000000101111000101000011111010000100;
	ram[149] = 82'b1010100100100001110011011111010111111011000011110111010000011000011011110010001000;
	ram[150] = 82'b1010100100001111010111000011110111011011100110001011110101011111011001001011000110;
	ram[151] = 82'b1010100011111100111100001000110100101000001101001011011000000111110111100110111000;
	ram[152] = 82'b1010100011101010100010101110000011000011000011101010001001111101100111011000000000;
	ram[153] = 82'b1010100011011000001010110011010100010011011110011011000111100010111101111110011001;
	ram[154] = 82'b1010100011000101110100011000011100000000101001000001000010010011111101110000000000;
	ram[155] = 82'b1010100010110011011111011101001101110100000100101011110110110111011011111000000000;
	ram[156] = 82'b1010100010100001001100000001011011011100101111011100011011001001111001000100110100;
	ram[157] = 82'b1010100010001110111010000100111000101001000111101010011101011000100011011000000000;
	ram[158] = 82'b1010100001111100101001100111011000100000011100000100110001101011000000111100010010;
	ram[159] = 82'b1010100001101010011010101000101110001100010111011111100001011000001101000000000000;
	ram[160] = 82'b1010100001011000001101001000101100111001000000001101100011111101100100000011100000;
	ram[161] = 82'b1010100001000110000001000111000111110100110111011001111011111000110001000000000000;
	ram[162] = 82'b1010100000110011110110100011110010010000111000100001010111100011011001111000101110;
	ram[163] = 82'b1010100000100001101101011110011110110111000000100110001100111010101101010111111011;
	ram[164] = 82'b1010100000001111100101110111000010001111110000110110101110000101011100110100000000;
	ram[165] = 82'b1010011111111101011111101101001110100000100001110110000101110101110100011010001000;
	ram[166] = 82'b1010011111101011011011000000110111101101001010110001011110001011011001000011110000;
	ram[167] = 82'b1010011111011001010111110001110001010010100010000110001110000001111011101111000000;
	ram[168] = 82'b1010011111000111010101111111101110101111110101000001011011001100010001000000000000;
	ram[169] = 82'b1010011110110101010101101010100011100110100110111001110110111000000110101000011000;
	ram[170] = 82'b1010011110100011010110110010000010110001101000100100110111111011100011100000010110;
	ram[171] = 82'b1010011110010001011001010110000000100000010101001111110101011110100001010110011000;
	ram[172] = 82'b1010011101111111011101010110010000011011001111111110101010011111100010000101010100;
	ram[173] = 82'b1010011101101101100010110010100110001101001111101010111110111101111100110001111000;
	ram[174] = 82'b1010011101011011101001101010110100111010011111001000011010010011110111110000000000;
	ram[175] = 82'b1010011101001001110001111110110000111011011111110010110001111000111100010111000000;
	ram[176] = 82'b1010011100110111111011101110001110000010000001100001000010111010100100101110000000;
	ram[177] = 82'b1010011100100110000110111000111111011001001100011001100011011011111100011010000011;
	ram[178] = 82'b1010011100010100010011011110111010001001001000011111000000111111101000011001001010;
	ram[179] = 82'b1010011100000010100001011111110000111000101000100100001001011010111101101001111000;
	ram[180] = 82'b1010011011110000110000111011010111100010100111001101100001111000010110011000100000;
	ram[181] = 82'b1010011011011111000001110001100010101100111110101110010001001110000001110001000000;
	ram[182] = 82'b1010011011001101010100000010000110010111000001111010011011100001110010110000000000;
	ram[183] = 82'b1010011010111011100111101100110110100010010001101111101111100000011111011000101000;
	ram[184] = 82'b1010011010101001111100110001100110101001110011011010110111000000000110111001001000;
	ram[185] = 82'b1010011010011000010011010000001010110011101001111010100001110001001101000100000011;
	ram[186] = 82'b1010011010000110101011001000011000011001010001100000101110110011010000000000000000;
	ram[187] = 82'b1010011001110101000100011010000010010011110010001010010110011100111111101000000000;
	ram[188] = 82'b1010011001100011011111000100111100101111110100101011101001000011010110011001110100;
	ram[189] = 82'b1010011001010001111011001000111100100100101100011010010110010000011010111000000000;
	ram[190] = 82'b1010011001000000011000100101110110000011010001111001111100100101010111100100000010;
	ram[191] = 82'b1010011000101110110111011011011100110110001100111101001100010011000010001100011111;
	ram[192] = 82'b1010011000011101010111101001100101010010110000100011101100111001100011101000000000;
	ram[193] = 82'b1010011000001011111001010000000101000001000111100011101101011111100001001101000000;
	ram[194] = 82'b1010010111111010011100001110101110100001101011111000110011001111001000100110110000;
	ram[195] = 82'b1010010111101001000000100101010111100000110111001000001101100010011001110011011000;
	ram[196] = 82'b1010010111010111100110010011110100011100011000110111101110010111000101100000000000;
	ram[197] = 82'b1010010111000110001101011001111001001011111000111101000010110111111110100110001101;
	ram[198] = 82'b1010010110110100110101110111011010111001100111110100110000100001100010001110000000;
	ram[199] = 82'b1010010110100011011111101100001101100001011111000101010000001111001001101111011000;
	ram[200] = 82'b1010010110010010001010111000000101101001101110110011100111110011010000011001011000;
	ram[201] = 82'b1010010110000000110111011010111000100010110010101010011010111111010101011010011000;
	ram[202] = 82'b1010010101101111100101010100011010001110111010100010010111010000100011001110000000;
	ram[203] = 82'b1010010101011110010100100100100000000010100111011110001000100000100101111001000000;
	ram[204] = 82'b1010010101001101000101001010111110000100010101101101010100100000110100101101010100;
	ram[205] = 82'b1010010100111011110111000111101001101100101001010001110000110010010010000011000000;
	ram[206] = 82'b1010010100101010101010011010010111000110001001010000001100011010101001101010000000;
	ram[207] = 82'b1010010100011001011111000010111011000101100001010111110010111110110111110100101001;
	ram[208] = 82'b1010010100001000010101000001001010100001011110111010011000111110101111101000010000;
	ram[209] = 82'b1010010011110111001100010100111010111010100110100111011001010011010011100100010101;
	ram[210] = 82'b1010010011100110000100111110000000100011101110110001001001011001000001110000000000;
	ram[211] = 82'b1010010011010100111110111100010001000001011001110001101100001001000110101001001111;
	ram[212] = 82'b1010010011000011111010001111100000101010100010100110101000011010100001011100100100;
	ram[213] = 82'b1010010010110010110110110111100100011111111001110111010010111101111010001000000000;
	ram[214] = 82'b1010010010100001110100110100010001100100001111000010111011000111010010101011010000;
	ram[215] = 82'b1010010010010000110100000101011101100011111001111111111101011000110110100100001000;
	ram[216] = 82'b1010010001111111110100101010111100111101111001110001110101101100111101000000011000;
	ram[217] = 82'b1010010001101110110110100100100100111010111000110101100100110010001001100100000111;
	ram[218] = 82'b1010010001011101111001110010001011001101000010001001101000110111001010100100000110;
	ram[219] = 82'b1010010001001100111110010011100100011001010010111111110111111010011010010100111000;
	ram[220] = 82'b1010010000111100000100001000100101000110101101110101101110010110100011110001011100;
	ram[221] = 82'b1010010000101011001011010001000100011100001100011111011111010100101111010110011101;
	ram[222] = 82'b1010010000011010010011101100110101110101101010110101101100110000010011110111010110;
	ram[223] = 82'b1010010000001001011101011011101111001110111011010001110110000010101100111011000000;
	ram[224] = 82'b1010001111111000101000011101100110100101100011011110000100000100101111100101100000;
	ram[225] = 82'b1010001111100111110100110010010000101010010000110101101100001010011100001110010001;
	ram[226] = 82'b1010001111010111000010011001100010110111000101110110011110011110111000110000000000;
	ram[227] = 82'b1010001111000110010001010011010010100111111110001101101111011001010000100011111000;
	ram[228] = 82'b1010001110110101100001011111010110000001111101010100011111111010110010111101100000;
	ram[229] = 82'b1010001110100100110010111101100001010110010000111010110001001110000110100010011000;
	ram[230] = 82'b1010001110010100000101101101101011010100111001010010100110000110000000000000000000;
	ram[231] = 82'b1010001110000011011001101111101000010010111011111111101001001100011011010110001000;
	ram[232] = 82'b1010001101110010101111000011001111000100000000010010010110110110110110000111000000;
	ram[233] = 82'b1010001101100010000101101000010100101000000110000001111001000000101011000010010001;
	ram[234] = 82'b1010001101010001011101011110101110101000001110001111011000110010101111011111100110;
	ram[235] = 82'b1010001101000000110110100110010010101111001111110011111101001101001101000000000000;
	ram[236] = 82'b1010001100110000010000111110110110101001110111000110010010010101110011101100000000;
	ram[237] = 82'b1010001100011111101100101000010000000110100101100000010011001011001010000101101111;
	ram[238] = 82'b1010001100001111001001100010010100110101110001000100110101111100100111000000100110;
	ram[239] = 82'b1010001011111110100111101100111010101001100100000101011011000110100010001111111000;
	ram[240] = 82'b1010001011101110000111000111110111010101111100100111111110110010101000111110000000;
	ram[241] = 82'b1010001011011101100111110011000001010111100001011010011001000010111011000111000000;
	ram[242] = 82'b1010001011001101001001101110001101011000001010110010101100111010000111000100010000;
	ram[243] = 82'b1010001010111100101100111001010001111000000110110011000001100101010100000100100001;
	ram[244] = 82'b1010001010101100010001010100000100110010011110101100110100100101100000000101001100;
	ram[245] = 82'b1010001010011011110110111110011100000100001101100011011101000000100000010101111000;
	ram[246] = 82'b1010001010001011011101111000001101101011111111110010001100010011010111010000000000;
	ram[247] = 82'b1010001001111011000110000001001111101010010010110010010001100110100111010001101011;
	ram[248] = 82'b1010001001101010101111011001011000000001010100100000111111100100001111101101011000;
	ram[249] = 82'b1010001001011010011010000000011100110101000011000101110100101111000000000000000000;
	ram[250] = 82'b1010001001001010000101110110010100001011001100011000100110011010101110011110110000;
	ram[251] = 82'b1010001000111001110010111010110100001011001101100111101110000101011111001110011101;
	ram[252] = 82'b1010001000101001100001001101110010111110010010111110011001010001000111110101110100;
	ram[253] = 82'b1010001000011001010000101111000110001000111010000010000110011111110011000110010111;
	ram[254] = 82'b1010001000001001000001011110100100011110001100111000010101101010101111110011010000;
	ram[255] = 82'b1010000111111000110011011100000100110010111100101011100001000110101000101000001101;
	ram[256] = 82'b1010000111101000100110100111011100001010010111111100001110100001101100000000000000;
	ram[257] = 82'b1010000111011000011011000000100001011100101011110010111011011110111001101000000000;
	ram[258] = 82'b1010000111001000010000100111001010111101010110010001110110100010000001001111011110;
	ram[259] = 82'b1010000110111000000111011011001110011011001111100111110110011010011000011111011000;
	ram[260] = 82'b1010000110100111111111011100100011011001110100010111011011001111101001111110111100;
	ram[261] = 82'b1010000110010111111000101010111111000101000011101100110110011010101110001000000000;
	ram[262] = 82'b1010000110000111110011000110011000011101011100101111111000110111101000011010000000;
	ram[263] = 82'b1010000101110111101110101110100101111110110111010010010010111000000001111010100101;
	ram[264] = 82'b1010000101100111101011100011011110000110110101010110011101001011001001100001101000;
	ram[265] = 82'b1010000101010111101001100100110110101110011100010000111010100000111011101110111011;
	ram[266] = 82'b1010000101000111101000110010100111100010110001010110110011011001111010101101011110;
	ram[267] = 82'b1010000100110111101001001100100101111010001000000101100101100110011011101000001101;
	ram[268] = 82'b1010000100100111101010110010101000011000101110001001101111001111110111001000110100;
	ram[269] = 82'b1010000100010111101101100100100110110000011000001101111111111110001100111011001101;
	ram[270] = 82'b1010000100000111110001100010010110011100011110101101001100010101111111100011010010;
	ram[271] = 82'b1010000011110111110110101011101110101100000011010111101110001001010010101000000000;
	ram[272] = 82'b1010000011100111111101000000100110001001101110010001001011010111101011110000000000;
	ram[273] = 82'b1010000011011000000100100000110010111011110111001000001101100111011010010111000000;
	ram[274] = 82'b1010000011001000001101001100001100010110001111001100011001110101101010101000111110;
	ram[275] = 82'b1010000010111000010111000010101001001000010010111011011011010111111100101110001111;
	ram[276] = 82'b1010000010101000100010000011111111011101010010101011010000101110111000010101101100;
	ram[277] = 82'b1010000010011000101110010000000110101101101100011011001110101000111001101111000000;
	ram[278] = 82'b1010000010001000111011100110110101101101101101110010010011101000001000101110000000;
	ram[279] = 82'b1010000001111001001010001000000010101101011100011010101001000110011100001000000000;
	ram[280] = 82'b1010000001101001011001110011100101001010000000000010001100000100111101001010101000;
	ram[281] = 82'b1010000001011001101010101001010011111100010100001001010111000101000111000000101001;
	ram[282] = 82'b1010000001001001111100101001000101011001010000101110101111011110100100010000010110;
	ram[283] = 82'b1010000000111010001111110010110001000010100011111100001010110101100001001000000000;
	ram[284] = 82'b1010000000101010100100000110001101110101110011111100100011000100111101011100000000;
	ram[285] = 82'b1010000000011010111001100011010010001100101000010110100001010011010110010111000000;
	ram[286] = 82'b1010000000001011010000001001110101101101010010001011011111011000111001101110000010;
	ram[287] = 82'b1001111111111011100111111001101110110100100001110011010001010100111001001011001000;
	ram[288] = 82'b1001111111101100000000110010110101001011101000100010111011111001000100000000000000;
	ram[289] = 82'b1001111111011100011010110100111111010010011101110101000001000100111001011101111000;
	ram[290] = 82'b1001111111001100110110000000000100110101010010010110001110001001100100000001111110;
	ram[291] = 82'b1001111110111101010010010011111100111100011001110000111001010000011010100001101001;
	ram[292] = 82'b1001111110101101101111110000011110001100010011101011110000110111000100001011001100;
	ram[293] = 82'b1001111110011110001110010101011111110000011010000000111101011110110001101100010011;
	ram[294] = 82'b1001111110001110101110000010111001011010110111110110100000110000000010000000010000;
	ram[295] = 82'b1001111101111111001110111000100010011010000001011011001110111000000000000000000000;
	ram[296] = 82'b1001111101101111110000110110010001011000011100010000111110011000001101101111000000;
	ram[297] = 82'b1001111101100000010011111011111110001100101011111010000001101111111101111100001111;
	ram[298] = 82'b1001111101010000111000001001011111100100010111011001000001010110011100100010000000;
	ram[299] = 82'b1001111101000001011101011110101100110011110011001011010011011111010001110010110111;
	ram[300] = 82'b1001111100110010000011111011011101110101111000010101001100011111010001101110101100;
	ram[301] = 82'b1001111100100010101011011111101010000001110001110000011001000000000000000000000000;
	ram[302] = 82'b1001111100010011010100001011001000001011000100101010001110010101010110011001001010;
	ram[303] = 82'b1001111100000011111101111101101111101011111011101110011011110101101110001100111000;
	ram[304] = 82'b1001111011110100101000110111011000100100111101011111000011101111000100110000000000;
	ram[305] = 82'b1001111011100101010100110111111001101110001010101110100000110101001011111101001000;
	ram[306] = 82'b1001111011010110000001111111001011001010111111000000110010101010000100110001010110;
	ram[307] = 82'b1001111011000110110000001101000011110110010110100001101000101010101000000000000000;
	ram[308] = 82'b1001111010110111011111100001011011010001101000001001000100000001110010100010110100;
	ram[309] = 82'b1001111010101000001111111100001001100100011100101010000001001100000110000100001001;
	ram[310] = 82'b1001111010011001000001011101000110010010111011011010111001100101110010011110000000;
	ram[311] = 82'b1001111010001001110100000100000111111001000001001111001010001111000001111000000000;
	ram[312] = 82'b1001111001111010100111110001000111000111010111000001010000011010110010101110001000;
	ram[313] = 82'b1001111001101011011100100011111011100110010011000111010001100000010101101010011001;
	ram[314] = 82'b1001111001011100010010011100011011110110001010101110110011100010101101010000000000;
	ram[315] = 82'b1001111001001101001001011010100000101011101001000000111100110110010110101111111000;
	ram[316] = 82'b1001111000111110000001011110000001110011010000011011110000100100101101000101100100;
	ram[317] = 82'b1001111000101110111010100110110101110001101011011101110100010011010011101110011101;
	ram[318] = 82'b1001111000011111110100110100110101011111100101010000000001010001100101101111010000;
	ram[319] = 82'b1001111000010000110000000111111000101101101001100001011100010010110111010000101000;
	ram[320] = 82'b1001111000000001101100011111110110000100110101011011001100101101011011100111000000;
	ram[321] = 82'b1001110111110010101001111100100110100001110001010101111011101111010001100011100011;
	ram[322] = 82'b1001110111100011101000011110000001111001001111011011100101011101000010001011110000;
	ram[323] = 82'b1001110111010100101000000011111110111000011101011011111001011000111101010101101000;
	ram[324] = 82'b1001110111000101101000101110010110011111111101101110000111111111001111100001100100;
	ram[325] = 82'b1001110110110110101010011101000000000100001100010101010101110000101001000000000000;
	ram[326] = 82'b1001110110100111101101001111110011011111011010110110001010100001010001010111100010;
	ram[327] = 82'b1001110110011000110001000110101001010001100111101011011011111000101010101010110111;
	ram[328] = 82'b1001110110001001110110000001011000110011010101010000110101101010001101001011011000;
	ram[329] = 82'b1001110101111010111011111111111010000010110101111100110110100101000111011011001001;
	ram[330] = 82'b1001110101101100000011000010000100111111110000110101110100000000011111111000001110;
	ram[331] = 82'b1001110101011101001011000111110001101011000001100001001110100101000111011110001011;
	ram[332] = 82'b1001110101001110010100010000111000101011000110101110110011000001010011100111100000;
	ram[333] = 82'b1001110100111111011110011101010001011111010010110100010111011110111011110101000011;
	ram[334] = 82'b1001110100110000101001101100110100001100011101111111000010101010000000000000000000;
	ram[335] = 82'b1001110100100001110101111111011000111000110011110110010001111000010011001001111011;
	ram[336] = 82'b1001110100010011000011010100111000001111111010110100111110100000110000101100010000;
	ram[337] = 82'b1001110100000100010001101101001001010010010100010100101000011010000000010100101000;
	ram[338] = 82'b1001110011110101100001001000000101010010010010001001101000110011000100111111010000;
	ram[339] = 82'b1001110011100110110001100101100011110111000011111010110101000101001101011001001000;
	ram[340] = 82'b1001110011011000000011000101011101001101010010111110001001011110001110100001100000;
	ram[341] = 82'b1001110011001001010101100111101001100010111010011110100011111010110011001010101000;
	ram[342] = 82'b1001110010111010101001001100000001000111000111001011101001100001001001010000110000;
	ram[343] = 82'b1001110010101011111101110010011100101110010011011000110100000101100010001110110011;
	ram[344] = 82'b1001110010011101010011011010110100000110001110110011011000001101100101011000000000;
	ram[345] = 82'b1001110010001110101010000100111110111110000001110001100111101000110100101000000000;
	ram[346] = 82'b1001110010000000000001110000110110110001101111000011111000100101101011100100010110;
	ram[347] = 82'b1001110001110001011010011110010011010010111101101110100110111001000000001001011000;
	ram[348] = 82'b1001110001100010110100001101001100111000011110111001100010000111111000101110111100;
	ram[349] = 82'b1001110001010100001110111101011011111010010011011100011100001101000000001111000000;
	ram[350] = 82'b1001110001000101101010101110111000110001101011101110111010101101001011100101011010;
	ram[351] = 82'b1001110000110111000111100001011011111001000111011000001001101000111000001010101000;
	ram[352] = 82'b1001110000101000100101010100111101101100010100111110101111101010011001010011100000;
	ram[353] = 82'b1001110000011010000100001001010111001011111101001110000101110011000011110100101111;
	ram[354] = 82'b1001110000001011100011111110011111101110110100000000111000101111100011100101110000;
	ram[355] = 82'b1001101111111101000100110100010000011000000000000010110100101101100111010000001011;
	ram[356] = 82'b1001101111101110100110101010100010001011101111110111101001101011110000011000011100;
	ram[357] = 82'b1001101111100000001001100001001100100100101011000101100101001010001100100011101000;
	ram[358] = 82'b1001101111010001101101011000001001001100111111101011000010010000000000000000000000;
	ram[359] = 82'b1001101111000011010010001111001111100001110110111000011111010000010000010011100101;
	ram[360] = 82'b1001101110110100111000000110011001001111110001111101011111011011101111111011101000;
	ram[361] = 82'b1001101110100110011110111101011101110110011010101101010000011001000001111101000000;
	ram[362] = 82'b1001101110011000000110110100010110100001001000011111110101101110111100000100001110;
	ram[363] = 82'b1001101110001001101111101010111100011100011001001111111010011100110110111110100111;
	ram[364] = 82'b1001101101111011011001100001000111001011100100100100010111000101000100101100000000;
	ram[365] = 82'b1001101101101101000100010110110000100000111000101000100000001110011100010110111000;
	ram[366] = 82'b1001101101011110110000001011110000000010001011011011110010000111100111010001110110;
	ram[367] = 82'b1001101101010000011100111111111111000000100110111001111101100011111101000000000000;
	ram[368] = 82'b1001101101000010001010110011010110001011000111010110001101101010110001010000010000;
	ram[369] = 82'b1001101100110011111001100101101110010001110011110011011011100101001111011110101000;
	ram[370] = 82'b1001101100100101101001010111000000000101111101110100011100010111100010010101000010;
	ram[371] = 82'b1001101100010111011010000111000100011010000001001100010000010011101111001111000000;
	ram[372] = 82'b1001101100001001001011110101110100000001100011101110010011100110011100001010011100;
	ram[373] = 82'b1001101011111010111110100011000111110001010100111110110000011100110101101111011000;
	ram[374] = 82'b1001101011101100110010001110111000011111001110000010110010100100001011111000101110;
	ram[375] = 82'b1001101011011110100110111000111110011111001010010110101110100011111110000000001111;
	ram[376] = 82'b1001101011010000011100100001010011101111100101011000101011100011000000000000000000;
	ram[377] = 82'b1001101011000010010011000111110000000011100110110011100110000000011110001001000000;
	ram[378] = 82'b1001101010110100001010101100001100111000110010101100100001011110110000001010000000;
	ram[379] = 82'b1001101010100110000011001110100011001010101110100011011011000000000000000000000000;
	ram[380] = 82'b1001101010010111111100101110101011110110000111111101110010001100110010100000000000;
	ram[381] = 82'b1001101010001001110111001100011111111000110100010111000110010100100110100111000000;
	ram[382] = 82'b1001101001111011110010100111111000010001110000110001010100100110011110100010000000;
	ram[383] = 82'b1001101001101101101111000000101101011110000111100011101000010001111001111011100111;
	ram[384] = 82'b1001101001011111101100010110111001100100111010101111001100000011010010110110000000;
	ram[385] = 82'b1001101001010001101010101010010100100010101010010010011001010110101001010010011000;
	ram[386] = 82'b1001101001000011101001111010110111111101101001111011010010111110011101000100001110;
	ram[387] = 82'b1001101000110101101010001000011100010111100101111011110111010110111000010101000111;
	ram[388] = 82'b1001101000100111101011010010111011111011101110011011100100100100110011101011100000;
	ram[389] = 82'b1001101000011001101101011010001110101011001001011000000100110000111000110101000000;
	ram[390] = 82'b1001101000001011110000011110001110010000011101010110010110101001100100011010010000;
	ram[391] = 82'b1001100111111101110100011110110011110100100010100101110011100010000010101111000000;
	ram[392] = 82'b1001100111101111111001011011111000100001010110100110100111111111111110100111000000;
	ram[393] = 82'b1001100111100001111111010101010100111111010001010100001011001110101110011110110101;
	ram[394] = 82'b1001100111010100000110001011000011011111110001110000000101110000101101110001000110;
	ram[395] = 82'b1001100111000110001101111100111100001010110000011100010110101101001110010000001000;
	ram[396] = 82'b1001100110111000010110101010111000001110100011001100111011000101100000010101100000;
	ram[397] = 82'b1001100110101010100000010100110001111111101101001100010101100011101011111100100101;
	ram[398] = 82'b1001100110011100101010111010100001101001011101010100010101011001001000110010000110;
	ram[399] = 82'b1001100110001110110110011100000000111111110111001010011111100101101000110000111011;
	ram[400] = 82'b1001100110000001000010111001001001010101011011110111001111100100010011011000010000;
	ram[401] = 82'b1001100101110011010000010001110011011011010001111011110101111011111110100000001000;
	ram[402] = 82'b1001100101100101011110100101111001001000100010100010001001010110101100010011011110;
	ram[403] = 82'b1001100101010111101101110101010011110010111000110000101100010000010100111000000000;
	ram[404] = 82'b1001100101001001111101111111111100110001000010001111001011000101100000100111000100;
	ram[405] = 82'b1001100100111100001111000101101100111000010111101100001000110010011000101111001011;
	ram[406] = 82'b1001100100101110100001000110011110000100000110110110101011111101100110111111011110;
	ram[407] = 82'b1001100100100000110100000010001001001011110000000001101101011010101010111000000000;
	ram[408] = 82'b1001100100010011000111111000101000101110110101100111101011110000000001111001000000;
	ram[409] = 82'b1001100100000101011100101001110100100010010110100001110011010011011010000101001000;
	ram[410] = 82'b1001100011110111110010010101100111101010000111011101011010110100011010010110001010;
	ram[411] = 82'b1001100011101010001000111011111010011111100001110110100001110110100110011011010111;
	ram[412] = 82'b1001100011011100100000011100100111000011110100110111000011111110010110100011001100;
	ram[413] = 82'b1001100011001110111000110111100110110110111110010111010100111101011011111100110101;
	ram[414] = 82'b1001100011000001010010001100110010110111110011010000000110111010011110100011110000;
	ram[415] = 82'b1001100010110011101100011100000100101000010111001010101111100111110100101000000000;
	ram[416] = 82'b1001100010100110000111100101010110101111111101010010011011111111011101000010100000;
	ram[417] = 82'b1001100010011000100011101000100001101110010101001111001011011100101110011101000111;
	ram[418] = 82'b1001100010001011000000100101011111101010100111101010100001011001111001010000100010;
	ram[419] = 82'b1001100001111101011110011100001001101000110010000000011011111000101001011000000000;
	ram[420] = 82'b1001100001101111111101001100011001110001111000110001111001010001010100010010101100;
	ram[421] = 82'b1001100001100010011100110110001001001011111011011001100011111111110010001010011111;
	ram[422] = 82'b1001100001010100111101011001010010000001111001111111110001101001101110000011101010;
	ram[423] = 82'b1001100001000111011110110101101101011011110100101110101001100011000000000000000000;
	ram[424] = 82'b1001100000111010000001001011010110001000100010010100111101110000100111001000000000;
	ram[425] = 82'b1001100000101100100100011010000100001110001011010011111100001111001111000000011000;
	ram[426] = 82'b1001100000011111001000100001110010111111011001101010010000100111101101101011001110;
	ram[427] = 82'b1001100000010001101101100010011010100100011011110101010110110000011010011010101000;
	ram[428] = 82'b1001100000000100010011011011110110010001101111000100111000001001000100001100000000;
	ram[429] = 82'b1001011111110110111010001101111110110011011010000010001010111010111000010100001011;
	ram[430] = 82'b1001011111101001100001111000101101111010010001100111110100010000100001001101100010;
	ram[431] = 82'b1001011111011100001010011011111101111001111000100000111110010011100100010111110101;
	ram[432] = 82'b1001011111001110110011110111101000100100111001100100110111110010100010011100010000;
	ram[433] = 82'b1001011111000001011110001011100111001101001111010100001010110000011011000000000000;
	ram[434] = 82'b1001011110110100001001010111110011100111100011000001011101010110011000100110010000;
	ram[435] = 82'b1001011110100110110101011100001000001011000101001101010010110000011111000000000000;
	ram[436] = 82'b1001011110011001100010011000011110101110010011111100000000001011101011111000100000;
	ram[437] = 82'b1001011110001100010000001100110000100111000001111010010010100000111001001101010101;
	ram[438] = 82'b1001011101111110111110111000110111101101101001111111011000001101001010001100011110;
	ram[439] = 82'b1001011101110001101110011100101110011101000111101110011101100100011011101110111011;
	ram[440] = 82'b1001011101100100011110111000001110101111101001001110101110111100100001101010111000;
	ram[441] = 82'b1001011101010111010000001011010001011101010100100010101000100011011000100011001011;
	ram[442] = 82'b1001011101001010000010010101110010000110111001000101111111001100101010000000000000;
	ram[443] = 82'b1001011100111100110101010111101001100110010100011011011010010010011100010011011000;
	ram[444] = 82'b1001011100101111101001010000110001111001100110100011000010110100011001001001111100;
	ram[445] = 82'b1001011100100010011110000001000101100001000101111011111111111011111100111011000000;
	ram[446] = 82'b1001011100010101010011101000011101111011001000111101111101010000100111011110000000;
	ram[447] = 82'b1001011100001000001010000110110101101001111000010010110000010111011101011000000000;
	ram[448] = 82'b1001011011111011000001011100000110001101100010001000010001111001001011111111000000;
	ram[449] = 82'b1001011011101101111001101000001001101000101010100010000101010101101101010101110111;
	ram[450] = 82'b1001011011100000110010101010111010100000000100001101110000001101000111100001000010;
	ram[451] = 82'b1001011011010011101100100100010010010110101111010110100111100111000101001000000000;
	ram[452] = 82'b1001011011000110100111010100001011110011001111011001101001111101100110110010001100;
	ram[453] = 82'b1001011010111001100010111010100000011010011010010010000111111100000011100111001111;
	ram[454] = 82'b1001011010101100011111010111001010010011010011111100010010100000001000110000000000;
	ram[455] = 82'b1001011010011111011100101010000100000111000111100010010010000100110111001100010111;
	ram[456] = 82'b1001011010010010011010110011000111111110100110011111011111000000111111011011000000;
	ram[457] = 82'b1001011010000101011001110010001111000001000101111000001100110110111100010000010001;
	ram[458] = 82'b1001011001111000011001100111010100011011100011110110011100110010011001110000000000;
	ram[459] = 82'b1001011001101011011010010010010010011001011011110011001000110110111110100011111001;
	ram[460] = 82'b1001011001011110011011110011000010000100110100100000011001110100010010000100000000;
	ram[461] = 82'b1001011001010001011110001001011110101101001100001001001101101110111101100011001101;
	ram[462] = 82'b1001011001000100100001010101100010100000100110011010101100100000100001011111110000;
	ram[463] = 82'b1001011000110111100101010111000111001100111100000010000101000001001000000000000000;
	ram[464] = 82'b1001011000101010101010001110000111000010000100010011111101000101011111110001110000;
	ram[465] = 82'b1001011000011101101111111010011100010000101101011111111111110110001100110110011011;
	ram[466] = 82'b1001011000010000110110011100000001101011011011000101110100001010000101100010111110;
	ram[467] = 82'b1001011000000011111101110010110001000011101000111011011000100111011111101000000000;
	ram[468] = 82'b1001010111110111000101111110100100101100101010011000000010100111010001010111100000;
	ram[469] = 82'b1001010111101010001110111111010111011011100011100100110101110110110111000000000000;
	ram[470] = 82'b1001010111011101011000110101000011000100011000011010011011011011110000001110111010;
	ram[471] = 82'b1001010111010000100011011111100001111100111111111100000001101001110110000001100101;
	ram[472] = 82'b1001010111000011101110111110101110111100111101001011001011110011010001111100001000;
	ram[473] = 82'b1001010110110110111011010010100011111010111010110100110001011010001110111000000000;
	ram[474] = 82'b1001010110101010001000011010111011001111010010001100011111010111111001110011010000;
	ram[475] = 82'b1001010110011101010110010111101111010011010010000000011001011111011111010110100011;
	ram[476] = 82'b1001010110010000100101001000111011000001101110111111100010100111010011110100000000;
	ram[477] = 82'b1001010110000011110100101110011000010100101111111100100101000110001110101111000000;
	ram[478] = 82'b1001010101110111000101001000000001101000000011111110011110111000111010100110101110;
	ram[479] = 82'b1001010101101010010110010101110001111000111011001010111100100101101101111011111000;
	ram[480] = 82'b1001010101011101101000010111100011000011111111110010100110101100100100000000000000;
	ram[481] = 82'b1001010101010000111011001101001111100111011111111010101111110001001111111111110011;
	ram[482] = 82'b1001010101000100001110110110110010000010011110000000001110111101000011101101100110;
	ram[483] = 82'b1001010100110111100011010100000100110100110000101110011111011111110111011000000000;
	ram[484] = 82'b1001010100101010111000100101000010111111101000001000011100010101110001000100100100;
	ram[485] = 82'b1001010100011110001110101001100110100011111011111001110101110011100011111011000011;
	ram[486] = 82'b1001010100010001100101100001101010000011111111011001101110011110111010101111110000;
	ram[487] = 82'b1001010100000100111101001101001000000010111001101000000110100010001100110010011000;
	ram[488] = 82'b1001010011111000010101101011111011100101000100101001101110101011110010110111000000;
	ram[489] = 82'b1001010011101011101110111101111110001110001110110000001101011001100001000000000000;
	ram[490] = 82'b1001010011011111001001000011001011100100110110111100001110110100001010110001110000;
	ram[491] = 82'b1001010011010010100011111011011101101110110010100010111010001001000001100111100011;
	ram[492] = 82'b1001010011000101111111100110101111110011100011100010111100111110100001100000000000;
	ram[493] = 82'b1001010010111001011100000100111011011010001111011101111110001001010101110111101001;
	ram[494] = 82'b1001010010101100111001010101111100001100010110010001101001010110001001011110010000;
	ram[495] = 82'b1001010010100000010111011001101100010010111110001101001001010010000001000111000000;
	ram[496] = 82'b1001010010010011110110010000000110011000011001111111010100101001001010001010010000;
	ram[497] = 82'b1001010010000111010101111001000101000111101110100011101011001010001011101010000111;
	ram[498] = 82'b1001010001111010110110010100100011001100110010111001100000010000010000000010000000;
	ram[499] = 82'b1001010001101110010111100010011011110100100000010010001101010010000011011100111111;
	ram[500] = 82'b1001010001100001111001100010101000101011110000000101100110111011011111100100000000;
	ram[501] = 82'b1001010001010101011100010101000101100001001101110101100101110010000001111010000011;
	ram[502] = 82'b1001010001001000111111111001101100100011100111100010110001001010010000000011111010;
	ram[503] = 82'b1001010000111100100100010000011000100010101100111011000000101111011000111111000000;
	ram[504] = 82'b1001010000110000001001011001000100001110111110111001100100101100111011101001000000;
	ram[505] = 82'b1001010000100011101111010011101010011001101111011110010101011100101000000111100101;
	ram[506] = 82'b1001010000010111010110000000000101110101000001100101000100000001010011011001001010;
	ram[507] = 82'b1001010000001010111101011110010001110011101110110100011100110100010010111111110011;
	ram[508] = 82'b1001001111111110100101101110001000001001001111001101011000101001000111000111100100;
	ram[509] = 82'b1001001111110010001110101111100100101010000001101110111001000111101101100110001101;
	ram[510] = 82'b1001001111100101111000100010100001101011000110001100100000111100001001110000000000;
	ram[511] = 82'b1001001111011001100011000110111001100010010010010101111110111011111110110100111011;
	ram[512] = 82'b1001001111001101001110011100101000000110001101111101101101111111110101000000000000;
	ram[513] = 82'b1001001111000000111010100011100111101110001101010010011101100111001011101111000000;
	ram[514] = 82'b1001001110110100100111011011110011010010010110000110101011001101110010010110101110;
	ram[515] = 82'b1001001110101000010101000101000110001011011000110000111100011001100100111100101000;
	ram[516] = 82'b1001001110011100000011011111011010010011000011011100101000110101101110010100101100;
	ram[517] = 82'b1001001110001111110010101010101011000011100110101001110010001101101000001010100001;
	ram[518] = 82'b1001001110000011100010100110110011011000000110000110110111011011001000101110000000;
	ram[519] = 82'b1001001101110111010011010011101110101100001010010010100110011101111110010000001001;
	ram[520] = 82'b1001001101101011000100110001010110111100101001000011001111111011100001000000000000;
	ram[521] = 82'b1001001101011110110110111111100111100110101001101001100111110111011111111010111000;
	ram[522] = 82'b1001001101010010101001111110011100000111111101100010101011011100000110000000000000;
	ram[523] = 82'b1001001101000110011101101101101110011111101110010001011001011010111000000000000000;
	ram[524] = 82'b1001001100111010010010001101011010101100111010011000010001100010011100000100000000;
	ram[525] = 82'b1001001100101110000111011101011010110000001101101001100111010100101111110100111000;
	ram[526] = 82'b1001001100100001111101011101101010101001111101110110000010000101011011000010000000;
	ram[527] = 82'b1001001100010101110100001110000100011100011000001110111011001111000000000000000000;
	ram[528] = 82'b1001001100001001101011101110100100001001001001011011110110110110000000000000000000;
	ram[529] = 82'b1001001011111101100011111111000011110011111111100011101001100111010001010101111000;
	ram[530] = 82'b1001001011110001011100111111011111011111111101100111010000100001101000110000000000;
	ram[531] = 82'b1001001011100101010110101111110001010010010001111111110100011011001001000000000000;
	ram[532] = 82'b1001001011011001010001001111110101001111010101100011101111000110000101010100000000;
	ram[533] = 82'b1001001011001101001100011111100101011101110110100001111001000001100000111001111000;
	ram[534] = 82'b1001001011000001001000011110111110000011100010111011110101001110001100000110000000;
	ram[535] = 82'b1001001010110101000101001101111001001000101000100000001001001000111001000000000000;
	ram[536] = 82'b1001001010101001000010101100010010110100001001101010110110101111011101000000000000;
	ram[537] = 82'b1001001010011101000000111010000101001111110011011010101110110010001101101100111000;
	ram[538] = 82'b1001001010010000111111110111001100000100011111010110000000011100011010110000011010;
	ram[539] = 82'b1001001010000100111111100011100010011100010011010010111101000010001101011100011011;
	ram[540] = 82'b1001001001111000111111111111000100000001011011111000011110011000011011111100001100;
	ram[541] = 82'b1001001001101101000001001001101011000000100001101001110001101000000100011001101011;
	ram[542] = 82'b1001001001100001000011000011010011000101001010100101010110010110110010110010010000;
	ram[543] = 82'b1001001001010101000101101011110111011100001101001100100100000011110001111001111000;
	ram[544] = 82'b1001001001001001001001000011010011010011001011110110110010011101111010001101100000;
	ram[545] = 82'b1001001000111101001101001001100001111000010100101001000100100110011101100001100001;
	ram[546] = 82'b1001001000110001010001111110011101111011001110110101110011111011100010011110001010;
	ram[547] = 82'b1001001000100101010111100010000011101010000110000001000000111100101001000010100111;
	ram[548] = 82'b1001001000011001011101110100001101110101110110101001111111000101001010100110100000;
	ram[549] = 82'b1001001000001101100100110100110111010000001110001010100011101010110000010010111001;
	ram[550] = 82'b1001001000000001101100100011111100001001010001110011000101000100000011111010000000;
	ram[551] = 82'b1001000111110101110101000001010110110100110111110000010011010101111101001001011111;
	ram[552] = 82'b1001000111101001111110001101000011000101001011001001111001101111010100101010111000;
	ram[553] = 82'b1001000111011110001000000110111100001101110011100101010100000001001100110100101000;
	ram[554] = 82'b1001000111010010010010101110111101100011000011001100101111000101000000000110110000;
	ram[555] = 82'b1001000111000110011110000101000010011001110110100110111010011010011101000001000101;
	ram[556] = 82'b1001000110111010101010001001000101101000101110111000100101010100001000001010100000;
	ram[557] = 82'b1001000110101110110110111011000011100100001010101011101001111001001100011100100101;
	ram[558] = 82'b1001000110100011000100011010110110100100111010010111010101010010110101010111110000;
	ram[559] = 82'b1001000110010111010010101000011011000000101011110110010111111001010100100001001001;
	ram[560] = 82'b1001000110001011100001100011101011010001101000101111001100111110100101111110000000;
	ram[561] = 82'b1001000101111111110001001100100011001111101101100001000010011010000001110000101000;
	ram[562] = 82'b1001000101110100000001100010111110010100011100111100110111110110000110000011011110;
	ram[563] = 82'b1001000101101000010010100110110111011011000110011001010001010100000001111111011000;
	ram[564] = 82'b1001000101011100100100011000001010111100011011000000110101110110111111110100010100;
	ram[565] = 82'b1001000101010000110110110110110011010110000000110110000111101000110111101001011000;
	ram[566] = 82'b1001000101000101001010000010101100100010111101001110101110001011000010000000000000;
	ram[567] = 82'b1001000100111001011101111011110010000000000001100110111001100100101011111110101001;
	ram[568] = 82'b1001000100101101110010100001111111001010101000010000100001100000000001010100101000;
	ram[569] = 82'b1001000100100010000111110101001111100000110100001010111111011001000111001101000000;
	ram[570] = 82'b1001000100010110011101110101011110000010011101000011010101001011100101111011101110;
	ram[571] = 82'b1001000100001010110100100010100110101101101110000000111101000110001000010011000101;
	ram[572] = 82'b1001000011111111001011111100100101000010100100001101111101100001100000000000000000;
	ram[573] = 82'b1001000011110011100100000011010100100001100101000011010001001000010001110100011000;
	ram[574] = 82'b1001000011100111111100110110110000101011111110000000100100001001001010001110101110;
	ram[575] = 82'b1001000011011100010110010110110100100100110110110001011101101110001011101010111000;
	ram[576] = 82'b1001000011010000110000100011011100001101011101110001101110011111001000000000000000;
	ram[577] = 82'b1001000011000101001011011100100011001000111000111101011010011100110111110100100011;
	ram[578] = 82'b1001000010111001100111000010000100111010110101111000110101011010000000101111100110;
	ram[579] = 82'b1001000010101110000011010011111101000111101001101000100011001111000110101000000000;
	ram[580] = 82'b1001000010100010100000010010000110110101101001011101111011010110110011100000101100;
	ram[581] = 82'b1001000010010110111101111100011110001001000011111110010000011101001010101111111111;
	ram[582] = 82'b1001000010001011011100010010111110101000000100111100110011011101101110000000000000;
	ram[583] = 82'b1001000001111111111011010101100011011010111011001111111111011011000011011100001101;
	ram[584] = 82'b1001000001110100011011000100001000100111100111100110000111100010011000100100011000;
	ram[585] = 82'b1001000001101000111011011110101001110110001011100001011100100110111101000000000000;
	ram[586] = 82'b1001000001011101011100100101000010101111001111001111110111010000111011111100010000;
	ram[587] = 82'b1001000001010001111110010111001110111100000001100010111101000010001001001000001011;
	ram[588] = 82'b1001000001000110100000110101001001100111111001111101001111110010000001101100100000;
	ram[589] = 82'b1001000000111011000011111110101110111011110101100001011100001001001001001000000000;
	ram[590] = 82'b1001000000101111100111110011111010100010110111000011011111010110110000000100100010;
	ram[591] = 82'b1001000000100100001100010100100111101010001101010110000000011000101100101111000000;
	ram[592] = 82'b1001000000011000110001100000110010011100100100110010111100001011001111000110000000;
	ram[593] = 82'b1001000000001101010111011000010110100110110011010001100001010111111011111011111101;
	ram[594] = 82'b1001000000000001111101111011001111010111111101010000000000110111100010010011010000;
	ram[595] = 82'b1000111111110110100101001001011001011010110100011100001010101000110011111010011001;
	ram[596] = 82'b1000111111101011001101000010101111100001010010111111101001100011111100000100100000;
	ram[597] = 82'b1000111111011111110101100111001101011010101010000111010010001000111100000000010011;
	ram[598] = 82'b1000111111010100011110110110101111110011010101000001110011100000110010000000000000;
	ram[599] = 82'b1000111111001001001000110001010001011111000110100110000010000001001010010100010001;
	ram[600] = 82'b1000111110111101110011010110101110001111000000011110000100010111111101101000000000;
	ram[601] = 82'b1000111110110010011110100111000010110001000111000010101000001100010111011100101101;
	ram[602] = 82'b1000111110100111001010100010001001111011000100011000000110010010110001100110000000;
	ram[603] = 82'b1000111110011011110111000111111111011111101001110001000000111111001011101011100011;
	ram[604] = 82'b1000111110010000100100011000100000001110100100000110010000110001100110111111100000;
	ram[605] = 82'b1000111110000101010010010011100110111111010011011101011011110101101001110000000101;
	ram[606] = 82'b1000111101111010000000111001001111100110010111111100110101110010111011011000010000;
	ram[607] = 82'b1000111101101110110000001001010110110101000110000000111110110111010111110100000001;
	ram[608] = 82'b1000111101100011100000000011110111100100110010110111011101111010010101110100000000;
	ram[609] = 82'b1000111101011000010000101000101101101011101100100101111001110110100011110111000011;
	ram[610] = 82'b1000111101001101000001110111110101111100101101111101001011001010000010011010000000;
	ram[611] = 82'b1000111101000001110011110001001011010011000000101100110011101110100001000001111001;
	ram[612] = 82'b1000111100110110100110010100101001100110100000000101011100000000000000000000000000;
	ram[613] = 82'b1000111100101011011001100010001101001101101011011100100101111111001110110001101000;
	ram[614] = 82'b1000111100100000001101011001110010000001100010101001111101001111000111101100100110;
	ram[615] = 82'b1000111100010101000001111011010011011101101010110100010111011000110010101000001000;
	ram[616] = 82'b1000111100001001110111000110101101111010001100001010011000110010111011000000000000;
	ram[617] = 82'b1000111011111110101100111011111101010001110001110110000111001111100000001100110111;
	ram[618] = 82'b1000111011110011100011011010111101000001101111100100110101011001110101101010000000;
	ram[619] = 82'b1000111011101000011010100011101001100011110101000000111000100111100011101011001000;
	ram[620] = 82'b1000111011011101010010010101111110110100010111101001101000011001100110101110111100;
	ram[621] = 82'b1000111011010010001010110001111000010010011001100101011010110010101010100111101000;
	ram[622] = 82'b1000111011000111000011110111010001111011011010100010011100011001111110101101100110;
	ram[623] = 82'b1000111010111011111101100110001000001011010010001110010111101100011101110100000011;
	ram[624] = 82'b1000111010110000110111111110010111000000100011100011000100101010011010110110000000;
	ram[625] = 82'b1000111010100101110010111111111010011010010011101011010101011110100101011111000000;
	ram[626] = 82'b1000111010011010101110101010101101111010011001101000000000000100000000100110000000;
	ram[627] = 82'b1000111010001111101010111110101101100001000100000100110010111100110111111001111000;
	ram[628] = 82'b1000111010000100100111111011110101101100110011010000100110001101101101001100100100;
	ram[629] = 82'b1000111001111001100101100010000010011110110111101111011010010100010001001100111001;
	ram[630] = 82'b1000111001101110100011110001001111011011010111011000101011111001101000101101010010;
	ram[631] = 82'b1000111001100011100010101001011001000010010110101101110000101000100010011100101000;
	ram[632] = 82'b1000111001011000100010001010011010111001000010100111001000101100010101110001001000;
	ram[633] = 82'b1000111001001101100010010100010001100000100001110111101001010000110000000011100101;
	ram[634] = 82'b1000111001000010100011000110111000111100110000001010011010100000100110000000000000;
	ram[635] = 82'b1000111000110111100100100010001100110100100100011011011101101100001100111000100011;
	ram[636] = 82'b1000111000101100100110100110001001001101000001111110010111100100100000000000000000;
	ram[637] = 82'b1000111000100001101001010010101010101001010010100000101011100000101100011001000000;
	ram[638] = 82'b1000111000010110101100100111101101001111011001100010001000110010010000011100000110;
	ram[639] = 82'b1000111000001011110000100101001100101000011001100110110001111100101111001011000000;
	ram[640] = 82'b1000111000000000110101001011000100111011011100100010011110101110000011011010000000;
	ram[641] = 82'b1000110111110101111010011001010011001011001110110010101000100111000001000111101000;
	ram[642] = 82'b1000110111101011000000001111110010000111011000101110011110000110011111101010010000;
	ram[643] = 82'b1000110111100000000110101110011110110011100111110111001011111001100000111101010101;
	ram[644] = 82'b1000110111010101001101110101010101011001001000100000100110111101111011100000100100;
	ram[645] = 82'b1000110111001010010101100100010001100100001011100100011011010000100001000010101101;
	ram[646] = 82'b1000110110111111011101111011001111111100011101011111011011010001101011010010010000;
	ram[647] = 82'b1000110110110100100110111010001100001111010011100100001110101110010000110010010111;
	ram[648] = 82'b1000110110101001110000100001000011000101011001100101000001101101000111000001001000;
	ram[649] = 82'b1000110110011110111010101111110000001101001000110110111101100010101100100011110111;
	ram[650] = 82'b1000110110010100000101100110010000010000001100001001010110101011100010110111010000;
	ram[651] = 82'b1000110110001001010001000100011110111110000000100000000111001110001010110111001001;
	ram[652] = 82'b1000110101111110011101001010011000100011111011011010101010011011001100001101100000;
	ram[653] = 82'b1000110101110011101001110111111001101101000101111111100010111101100011110010011000;
	ram[654] = 82'b1000110101101000110111001100111110100111110011100000100010001110000010010101000010;
	ram[655] = 82'b1000110101011110000101001001100011000101100110010111110001111001000111010111001000;
	ram[656] = 82'b1000110101010011010011101101100011110011000100111000001110110011110000000010000000;
	ram[657] = 82'b1000110101001000100010111000111100000101100110001011111101100000100101001110111101;
	ram[658] = 82'b1000110100111101110010101011101001100101001100001011000010011000000010001010000000;
	ram[659] = 82'b1000110100110011000011000101100111101000001110010110011101000011101011001101100011;
	ram[660] = 82'b1000110100101000010100000110110010100000000011100011000000001101110010011100000000;
	ram[661] = 82'b1000110100011101100101101111000110111011101011101110011011110011111110100101000000;
	ram[662] = 82'b1000110100010010110111111110100000110000010000110101011110011001010010010101110000;
	ram[663] = 82'b1000110100001000001010110100111100101101101111110000000100010001011100110010000011;
	ram[664] = 82'b1000110011111101011110010010010110101010010011110011011010000001001010011101000000;
	ram[665] = 82'b1000110011110010110010010110101010111001110001001011000110110010100001011010001101;
	ram[666] = 82'b1000110011101000000111000001110110001101011111101001110001100000010001100100101010;
	ram[667] = 82'b1000110011011101011100010011110100011101001011011100100111000001011001101100111001;
	ram[668] = 82'b1000110011010010110010001100100010011011001000111000011110111011111101100101100000;
	ram[669] = 82'b1000110011001000001000101011111100000000000100010001011110111001110010110110110011;
	ram[670] = 82'b1000110010111101011111110001111101111111001101101101011111000110011010011110111110;
	ram[671] = 82'b1000110010110010110111011110100100010010010001101101101011110110010001111001001111;
	ram[672] = 82'b1000110010101000001111110001101011010000011101111001100101101000111011011101100000;
	ram[673] = 82'b1000110010011101101000101011001111101110011011010111001001000011111011110001101000;
	ram[674] = 82'b1000110010010011000010001011001101100111010110000010011101101111000110010010010110;
	ram[675] = 82'b1000110010001000011100010001100001110000110010000101001010010011001010000101111011;
	ram[676] = 82'b1000110001111101110110111110001000000110111010101101001000100010011000110111110100;
	ram[677] = 82'b1000110001110011010010010000111101000011010110010100011100001111110100011101011011;
	ram[678] = 82'b1000110001101000101110001001111101011101000000110111101010010110001100011101010000;
	ram[679] = 82'b1000110001011110001010101001000101010001100011110100110000110110100101010100010101;
	ram[680] = 82'b1000110001010011100111101110010001011000110101001111011110101101110101101100001000;
	ram[681] = 82'b1000110001001001000101011001011101010100101001001111001011001011101010000011111000;
	ram[682] = 82'b1000110000111110100011101010100110110111011000111110110010101000100000010110001110;
	ram[683] = 82'b1000110000110100000010100001101001000111000011010010111110101000010010100001001101;
	ram[684] = 82'b1000110000101001100001111110100001011010000101111111011100100111000110100000000000;
	ram[685] = 82'b1000110000011111000010000001001100001101110100011100101000001010010010001100111000;
	ram[686] = 82'b1000110000010100100010101001100101000110100010100010011100110111111110000000111010;
	ram[687] = 82'b1000110000001010000011110111101001011100000000100000100101111010011110100101111011;
	ram[688] = 82'b1000101111111111100101101011010101101100111010101111100001011100000100110000000000;
	ram[689] = 82'b1000101111110101001000000100100101111011101111001100011110100110101001100100111001;
	ram[690] = 82'b1000101111101010101011000011010110101000001000011111111000100001110010000110000000;
	ram[691] = 82'b1000101111100000001110100111100100010010001110000101110001000001001101000000011111;
	ram[692] = 82'b1000101111010101110010110001001011110111001100110110011101111000111010010001011100;
	ram[693] = 82'b1000101111001011010111100000001001011011011100011101110000001010001011011010110011;
	ram[694] = 82'b1000101111000000111100110100011001100000011011110001111110000001000011011100110110;
	ram[695] = 82'b1000101110110110100010101101111001000100101100000101010110110110011101011000000000;
	ram[696] = 82'b1000101110101100001001001100100100001101111110110100010101001000111101000100011000;
	ram[697] = 82'b1000101110100001110000010000010111111011101100101001001001111001000100001000010111;
	ram[698] = 82'b1000101110010111010111111001001111111000000001010110011100000010100010000000000000;
	ram[699] = 82'b1000101110001101000000000111001001011111110000101011001010101010001110110011101000;
	ram[700] = 82'b1000101110000010101000111010000001010111000011010001011110110001010100111101011100;
	ram[701] = 82'b1000101101111000010010010001110011001001100000111011111010011111110110111100001111;
	ram[702] = 82'b1000101101101101111100001110011100010101001100110101001001110101000011000110110000;
	ram[703] = 82'b1000101101100011100110101111111001000011001000001110100010011110000011101110010001;
	ram[704] = 82'b1000101101011001010001110110000110010101101100100001100000110010010111111011000000;
	ram[705] = 82'b1000101101001110111101100001000000010110110101010110011101010111100100000001010001;
	ram[706] = 82'b1000101101000100101001110000100011101101011000110010011111101001010001110000111110;
	ram[707] = 82'b1000101100111010010110100100101101000000101000101010011110000010101000001010011001;
	ram[708] = 82'b1000101100110000000011111101011001010100101010100010111001010100010010110100000000;
	ram[709] = 82'b1000101100100101110001111010100100110101001110101100010011101100001011001101101111;
	ram[710] = 82'b1000101100011011100000011100001100001010111010111100111011110111110000000000000000;
	ram[711] = 82'b1000101100010001001111100010001100011011000101001011100111111101110100001110111000;
	ram[712] = 82'b1000101100000110111111001100100001110010110100010011100111111101100110001001000000;
	ram[713] = 82'b1000101011111100101111011011001000111100000001100100000101111110011000000000000000;
	ram[714] = 82'b1000101011110010100000001101111110100001000001011110110100100101011101100110000000;
	ram[715] = 82'b1000101011101000010001100100111111001100100011110100011001100100110110011010001000;
	ram[716] = 82'b1000101011011110000011100000001000000110000011100010110100110111001111000010111100;
	ram[717] = 82'b1000101011010011110101111111010101011100110110001011100010101101010101100101101000;
	ram[718] = 82'b1000101011001001101001000010100100011001001010111111111100110011111100000110000000;
	ram[719] = 82'b1000101010111111011100101001110000101111000100100110000001010101111001011100110011;
	ram[720] = 82'b1000101010110101010000110100111000000011110100010100000110010100100000101011110000;
	ram[721] = 82'b1000101010101011000101100011110110101000100000111010000010000100110110011100101111;
	ram[722] = 82'b1000101010100000111010110110101001001010111001000010011000110101011100011011000010;
	ram[723] = 82'b1000101010010110110000101101001100110101001110011011001001010111100111000000000000;
	ram[724] = 82'b1000101010001100100111000111011101111001111011011011110001101000111110110111000100;
	ram[725] = 82'b1000101010000010011110000101011001000111111111101010101010111001010100111000000000;
	ram[726] = 82'b1000101001111000010101100110111011001110110101001111111101011010100011100011000110;
	ram[727] = 82'b1000101001101110001101101100000000111110010000110001101110100110001100101000000000;
	ram[728] = 82'b1000101001100100000110010100100111100010100100011110100011010011100100111000000000;
	ram[729] = 82'b1000101001011001111111100000101011010000010101011011101101011101011000100111111000;
	ram[730] = 82'b1000101001001111111001010000001000111000101000001011000110111001111110111011110000;
	ram[731] = 82'b1000101001000101110011100010111101001100111011011100011101111110010011110101000000;
	ram[732] = 82'b1000101000111011101110011001000101011011000110110111001110010001100110011101100100;
	ram[733] = 82'b1000101000110001101001110010011101011101011111111011111110101010101011000001111101;
	ram[734] = 82'b1000101000100111100101101111000010111110110000001111000111111010010010000000000000;
	ram[735] = 82'b1000101000011101100010001110110010010110000000111000111101010011100100101111111011;
	ram[736] = 82'b1000101000010011011111010001101000110010101110001100000011011000110010011000100000;
	ram[737] = 82'b1000101000001001011100110111100010010000111110010001101100101111001001000000000000;
	ram[738] = 82'b1000100111111111011011000000011100011100111010011000011111101011010110110000110000;
	ram[739] = 82'b1000100111110101011001101100010011101111010111110110101000000110000110111011111000;
	ram[740] = 82'b1000100111101011011000111011000100111101100000001110111011011110101111111100000000;
	ram[741] = 82'b1000100111100001011000101100101100111100110110101010100011111110011111110011000000;
	ram[742] = 82'b1000100111010111011001000001001000100011010111110101010010100010010000101011110000;
	ram[743] = 82'b1000100111001101011001111000010101000011001101011011010010110101001110010000011011;
	ram[744] = 82'b1000100111000011011011010010001110011011011111111101100100001010111010000010011000;
	ram[745] = 82'b1000100110111001011101001110110010011010111110011111000100001001111011111010011000;
	ram[746] = 82'b1000100110101111011111101101111101011101011000011010111011011111111000110010111110;
	ram[747] = 82'b1000100110100101100010101111101100011010101001111100110111001011010100010001101000;
	ram[748] = 82'b1000100110011011100110010011111100100110110111000111011010000111010101111010100000;
	ram[749] = 82'b1000100110010001101010011010101010000011010000101110011110010111000010010010110001;
	ram[750] = 82'b1000100110000111101111000011110010100000011010011001011111000010010000001110011110;
	ram[751] = 82'b1000100101111101110100001111010010011100000110100111011101000001110111000011010101;
	ram[752] = 82'b1000100101110011111001111101000110110000001111011110011110010101110110000111010000;
	ram[753] = 82'b1000100101101010000000001101001100010111000111111100100011101101100001110111000001;
	ram[754] = 82'b1000100101100000000110111111100000001011011011110011111101111100001111010100001010;
	ram[755] = 82'b1000100101010110001110010011111111001000001111100111100011011110000000001011000101;
	ram[756] = 82'b1000100101001100010110001010100110100100100111010010001111111001111010110011100000;
	ram[757] = 82'b1000100101000010011110100011010010100101001011001101101000101010011010001001000000;
	ram[758] = 82'b1000100100111000100111011110000000111101010110000010101010010101110110010110101010;
	ram[759] = 82'b1000100100101110110000111010101110001110001000100111111110110111001011011000000000;
	ram[760] = 82'b1000100100100100111010111001010111010100100010111100101101001110101111100100001000;
	ram[761] = 82'b1000100100011011000101011001111001001101111101011001100110111101011011100101000000;
	ram[762] = 82'b1000100100010001010000011100010000111000001000101101011111011101010110001110110110;
	ram[763] = 82'b1000100100000111011100000000011011010001001101111001100011101010010110101000000000;
	ram[764] = 82'b1000100011111101101000000110010101110011001101010001000100010110100010100010100000;
	ram[765] = 82'b1000100011110011110100101101111100100110000001111000111101111111100111101110011111;
	ram[766] = 82'b1000100011101010000001110111001101011111111010000011100110111111001011111111110110;
	ram[767] = 82'b1000100011100000001111100010000101000101000000101111000111011101000111001110100011;
	ram[768] = 82'b1000100011010110011101101110100000010101010111111100001011111011110100010100000000;
	ram[769] = 82'b1000100011001100101100011100011100010001011001100111001100000111110010011010001111;
	ram[770] = 82'b1000100011000010111011101011110101111001110111100100100100010010111010100010100010;
	ram[771] = 82'b1000100010111001001011011100101010001111111011011101001110111111100001000100110011;
	ram[772] = 82'b1000100010101111011011101110110110010101000110101010111110111011000001111000111100;
	ram[773] = 82'b1000100010100101101100100010010111001011010010010100111001001000010101111011011111;
	ram[774] = 82'b1000100010011011111101110111001001110100101111001011101111011001110000111110101110;
	ram[775] = 82'b1000100010010010001111101101001011101111011001110010000001000100010110000001000000;
	ram[776] = 82'b1000100010001000100010000100011001000111101001010111100101110011100100011001000000;
	ram[777] = 82'b1000100001111110110100111100101111110111011100001100011010111100111100000101100101;
	ram[778] = 82'b1000100001110101001000010110001100001011111100010111101011111000000101010100000110;
	ram[779] = 82'b1000100001101011011100010000101011111111110011010110111110011011000000101011001000;
	ram[780] = 82'b1000100001100001110000101100001011111100001100100111011100001011101001101010000100;
	ram[781] = 82'b1000100001011000000101101000101001000101111101001001001001000100000010110010011000;
	ram[782] = 82'b1000100001001110011011000110000000100010010001001000010001000101101100101110000010;
	ram[783] = 82'b1000100001000100110001000100001110111011011111111001011110010100011100111011000001;
	ram[784] = 82'b1000100000111011000111100011010010001101111100110111100001010111111001010000000000;
	ram[785] = 82'b1000100000110001011110100011000111000100101100011000100000011101011101101010110111;
	ram[786] = 82'b1000100000100111110110000011101011000001100000000000011000110000001101101110111110;
	ram[787] = 82'b1000100000011110001110000100111010010101000011111001011100011100011011100001001000;
	ram[788] = 82'b1000100000010100100110100110110010100001111000010001000011100010011110100001011100;
	ram[789] = 82'b1000100000001010111111101001010000101111101010000101000010110000101001001000011000;
	ram[790] = 82'b1000100000000001011001001100010010000110011101000011000010111100000111100100111010;
	ram[791] = 82'b1000011111110111110011001111110011101110101011100100111111100101111100101101001000;
	ram[792] = 82'b1000011111101110001101110011110011001100001010010010011010000010011110101011000000;
	ram[793] = 82'b1000011111100100101000111000001100110001111001000110100011001001101011110110010101;
	ram[794] = 82'b1000011111011011000100011100111110000100011010010101000011111010101001010001110000;
	ram[795] = 82'b1000011111010001100000100010000100101000100011001100101101001000110111101011000000;
	ram[796] = 82'b1000011111000111111101000111011100110010011101000100000110101010000011111101011100;
	ram[797] = 82'b1000011110111110011010001101000100000111101010011010111110111110110111001011000000;
	ram[798] = 82'b1000011110110100110111110010111000001110000000110101100111101111111011001110000000;
	ram[799] = 82'b1000011110101011010101111000110101011010110010001000101001100000100010101100001101;
	ram[800] = 82'b1000011110100001110100011110111001010100100000110000011101101011100000000000000000;
	ram[801] = 82'b1000011110011000010011100101000001100010000010001110011111110110110000110001001000;
	ram[802] = 82'b1000011110001110110011001011001010011001110000000101100111000000100110110100110110;
	ram[803] = 82'b1000011110000101010011010001010001111110000101011000110110111011000000010100010011;
	ram[804] = 82'b1000011101111011110011110111010100100110001100000111101111000111111000001111100000;
	ram[805] = 82'b1000011101110010010100111101001111111010010000000001001100011111111000110111111101;
	ram[806] = 82'b1000011101101000110110100011000001100010101111100110001011111000111001100011100110;
	ram[807] = 82'b1000011101011111011000101000100101110111111011110010111000001111111100101000000000;
	ram[808] = 82'b1000011101010101111011001101111010100010111111001001010111111000100010010001001000;
	ram[809] = 82'b1000011101001100011110010010111101001101010110100110100000111101100000111110010111;
	ram[810] = 82'b1000011101000011000001110111101010010000011001110111010111101000111110000000000000;
	ram[811] = 82'b1000011100111001100101111011111111010110010001101001100001010001111010111111110101;
	ram[812] = 82'b1000011100110000001010011111111001101110101000010000001110110001101000100100000000;
	ram[813] = 82'b1000011100100110101111100011010111000100001101001001111110101111110000000000111000;
	ram[814] = 82'b1000011100011101010101000110010011110001110101100010101111000101101010101010010010;
	ram[815] = 82'b1000011100010011111011001000101101100010111100010111011000010000101000111010101000;
	ram[816] = 82'b1000011100001010100001101010100001101000100001100101010001100110011110000010010000;
	ram[817] = 82'b1000011100000001001000101011101101010011111010011011110011001000110111111100111000;
	ram[818] = 82'b1000011011110111110000001100001101110110110001011000111010100000000100011101101110;
	ram[819] = 82'b1000011011101110011000001100000000100011000110000101110000000100000110101110101000;
	ram[820] = 82'b1000011011100101000000101011000010101011001101010011001100010100111011110011011100;
	ram[821] = 82'b1000011011011011101001101001010001100001110000110110011101100001001101000010111000;
	ram[822] = 82'b1000011011010010010011000110101010011001101111100101101101011011101111000110001010;
	ram[823] = 82'b1000011011001000111101000011001010001011110111010000010111100101111100001100100001;
	ram[824] = 82'b1000011010111111100111011110101111000000111110000011101100000110010011101000000000;
	ram[825] = 82'b1000011010110110010010011001010101110010011010001110100110010100110010011011100111;
	ram[826] = 82'b1000011010101100111101110010111011011001111010111111101000000000011110111011011010;
	ram[827] = 82'b1000011010100011101001101011011110000001001111011010011011000000000000000000000000;
	ram[828] = 82'b1000011010011010010110000010111010001000001101011010010001101000101001111100100000;
	ram[829] = 82'b1000011010010001000010111001001101011110101000111010001011000101100000011000001000;
	ram[830] = 82'b1000011010000111110000001110010101110100100111100101000011010010101110110001001010;
	ram[831] = 82'b1000011001111110011110000010001111101011000010001001000111101010100111000100101101;
	ram[832] = 82'b1000011001110101001100010100111000110010100111110101010000111111011000101101000000;
	ram[833] = 82'b1000011001101011111011000110001110100001111011100001011100011101110010000101001101;
	ram[834] = 82'b1000011001100010101010010110001110001111110100011110111000100110000110000100001110;
	ram[835] = 82'b1000011001011001011010000100110101010011011110010100101101111011000001101101110101;
	ram[836] = 82'b1000011001010000001010010010000001000100011000111100100111111110111101111101110100;
	ram[837] = 82'b1000011001000110111010111101101110011111111111000100001010101101100101110101101000;
	ram[838] = 82'b1000011000111101101100000111111011110011001101010110010101000101011001010010000000;
	ram[839] = 82'b1000011000110100011101110000100101100001101101101111101011110011110111101101001011;
	ram[840] = 82'b1000011000101011001111110111101001111001000010000001110001010001011011001011011000;
	ram[841] = 82'b1000011000100010000010011101000101011101011111111100110001111001000001000000000000;
	ram[842] = 82'b1000011000011000110101100000110110000010111000001111000100101100010001100101001110;
	ram[843] = 82'b1000011000001111101001000010111001000010110111110100011111111000101001010111000000;
	ram[844] = 82'b1000011000000110011101000011001011110111011111100001101001110111100000110110000100;
	ram[845] = 82'b1000010111111101010001100001101011111011000100000000100100001000101001000000000000;
	ram[846] = 82'b1000010111110100000110011110010110101000001101101101010110011010110111101111101010;
	ram[847] = 82'b1000010111101010111011111001001001011001111000110010111010000011000011010111000000;
	ram[848] = 82'b1000010111100001110001110010000001010001000110000110011001100101001001110000000000;
	ram[849] = 82'b1000010111011000101000001000111100000011101010010010001001001100111010001111001000;
	ram[850] = 82'b1000010111001111011110111101110111100111101011000010110110001011111100111101101010;
	ram[851] = 82'b1000010111000110010110010000110000100100110110100100011110111010011011010011100101;
	ram[852] = 82'b1000010110111101001110000001100100110001111010001000000100100010110001110001001100;
	ram[853] = 82'b1000010110110100000110010000010001101011100111110000101110101011111001010010010001;
	ram[854] = 82'b1000010110101010111110111100110100010100111010110110100010000011101010101100110000;
	ram[855] = 82'b1000010110100001111000000111001010111111100001110001100100011001011101110101000000;
	ram[856] = 82'b1000010110011000110001101111010010010100110100111011010100101110001100001111111000;
	ram[857] = 82'b1000010110001111101011110101001000100111000110000101010011010000011001101000101011;
	ram[858] = 82'b1000010110000110100110011000101010100000010111111111110010111011100110000000000000;
	ram[859] = 82'b1000010101111101100001011001110101111001011001001011110110011010000111010110011001;
	ram[860] = 82'b1000010101110100011100111000101000010001000010111101011100111110011111101100000000;
	ram[861] = 82'b1000010101101011011000110100111110101100011101110101110111000100001110010101000000;
	ram[862] = 82'b1000010101100010010101001110110111011111010010011000010110110000011010101000111110;
	ram[863] = 82'b1000010101011001010010000110001111010101001011110000000111100111000110000100111011;
	ram[864] = 82'b1000010101010000001111011011000100001000010011101001000010100011010110100110100000;
	ram[865] = 82'b1000010101000111001101001101010011110011000011010101101100001100100000011010111000;
	ram[866] = 82'b1000010100111110001011011100111010101000000100100101100111000000100001010110111010;
	ram[867] = 82'b1000010100110101001010001001110111010110010111011001011100111100100010011010111011;
	ram[868] = 82'b1000010100101100001001010100000111000101001100001000010101001010110111000010101100;
	ram[869] = 82'b1000010100100011001000111011100110111100001001111101000010010001000100000011000000;
	ram[870] = 82'b1000010100011010001001000000010100110111000110000101010110001111011110001111110010;
	ram[871] = 82'b1000010100010001001001100010001110011000001010000001010011110001101100101000000000;
	ram[872] = 82'b1000010100001000001010100001010001000001110001110001100010101000100100110101111000;
	ram[873] = 82'b1000010011111111001011111101011010010110101011110100000000011101101000000011000000;
	ram[874] = 82'b1000010011110110001101110110100111100000000000100111111000100100001001001010000000;
	ram[875] = 82'b1000010011101101010000001100110110110100110110000110110110110000011110001011100011;
	ram[876] = 82'b1000010011100100010011000000000101000101000010000001001100110110100101111001011100;
	ram[877] = 82'b1000010011011011010110010000010000001110010101010111111011100110111100010001110011;
	ram[878] = 82'b1000010011010010011001111101010101011011000110000100000011011010101110000000000000;
	ram[879] = 82'b1000010011001001011110000111010011000011011100100100111011100000001100000010001000;
	ram[880] = 82'b1000010011000000100010101110000101111000011110110100110100100101100011000101010000;
	ram[881] = 82'b1000010010110111100111110001101011111001000011110110000111011010100110010100011000;
	ram[882] = 82'b1000010010101110101101010010000010101010011111110000001010101110011110011100001110;
	ram[883] = 82'b1000010010100101110011001111000111110010011000101001010110001011101010101110001000;
	ram[884] = 82'b1000010010011100111001101000111000011100110110101001000011010000100110111100000000;
	ram[885] = 82'b1000010010010100000000011111010011000011100101011000001111110111100101001100011011;
	ram[886] = 82'b1000010010001011000111110010010100011001100001110100111100000000100000101000010110;
	ram[887] = 82'b1000010010000010001111100001111010011111001010011000001000100101101010000101100111;
	ram[888] = 82'b1000010001111001010111101110000010100001110010111011111101011011111000000000000000;
	ram[889] = 82'b1000010001110000100000010110101010111100000111101111100011100011100011101011000000;
	ram[890] = 82'b1000010001100111101001011011110000100010010100100111110001111101011111011011110110;
	ram[891] = 82'b1000010001011110110010111101010001010101111100000010000111010110111000000000000000;
	ram[892] = 82'b1000010001010101111100111011001010111111000101101100001000001011010110000111100100;
	ram[893] = 82'b1000010001001101000111010101011010101100100010111100011101000010101101000010000001;
	ram[894] = 82'b1000010001000100010010001011111110111010010000000111101001101111110000000000000000;
	ram[895] = 82'b1000010000111011011101011110110100011101111010101011110000001100011111101010111000;
	ram[896] = 82'b1000010000110010101001001101111001000000110011011100100110001000110010101010000000;
	ram[897] = 82'b1000010000101001110101011001001010111111100110110101011110111010000000001000110001;
	ram[898] = 82'b1000010000100001000010000000100111010000111011100010001011101100110010010011110000;
	ram[899] = 82'b1000010000011000001111000100001011111000011010100001001110000100100101111100101011;
	ram[900] = 82'b1000010000001111011100100011110110100000011000011001011110101001000110000100100000;
	ram[901] = 82'b1000010000000110101010011111100100110011011010111011011000111000110100011100001101;
	ram[902] = 82'b1000001111111101111000110111010100000010111000101101101011011100100010110101111010;
	ram[903] = 82'b1000001111110101000111101011000010010011011100110000010101111001111001110101111101;
	ram[904] = 82'b1000001111101100010110111010101101010000100001000100100011100101111110110101101000;
	ram[905] = 82'b1000001111100011100110100110010010100101110000101001011000111100111101100000100101;
	ram[906] = 82'b1000001111011010110110101101101111100101101010101011100010101110011011001010000000;
	ram[907] = 82'b1000001111010010000111010001000010010101111011100100111001001000000011000111001011;
	ram[908] = 82'b1000001111001001011000010000001000100011000010000100111110011010101101110100000000;
	ram[909] = 82'b1000001111000000101001101010111111111001101101101101100111001000100010111000101001;
	ram[910] = 82'b1000001110110111111011100001100101101101100101110101100000100011000010101101100110;
	ram[911] = 82'b1000001110101111001101110011111000000101010111011011011111011010001010001110110101;
	ram[912] = 82'b1000001110100110100000100001110100101110100101010001101100001110101010000011110000;
	ram[913] = 82'b1000001110011101110011101011011000111101101100000101000000100101000000110001101000;
	ram[914] = 82'b1000001110010101000111010000100010111010001001000100010000010110010011100100110110;
	ram[915] = 82'b1000001110001100011011010001010000010010010001111010011111011010001101010110111000;
	ram[916] = 82'b1000001110000011101111101101011110110100101100110001000101011011000110100100001100;
	ram[917] = 82'b1000001101111011000100100101001011110110111100110010001010110011010011100101110111;
	ram[918] = 82'b1000001101110010011001111000010101100001011111010011001000010001100000010000001110;
	ram[919] = 82'b1000001101101001101111100110111001100011101100110110010101000101010111001000001011;
	ram[920] = 82'b1000001101100001000101110000110101010011111100111010111111110011001011101000000000;
	ram[921] = 82'b1000001101011000011100010110000111010100101101010011100111110000111000000000000000;
	ram[922] = 82'b1000001101001111110011010110101100100011100110000001000001010000011000010000111110;
	ram[923] = 82'b1000001101000111001010110010100010110001000100110000100101110011011001110011001111;
	ram[924] = 82'b1000001100111110100010101001101000000111000100111111111101011000101000001000101100;
	ram[925] = 82'b1000001100110101111010111011111010010110100010111101101001010001011010100100101111;
	ram[926] = 82'b1000001100101101010011101001010111010000101010111010010011010011110000111001100010;
	ram[927] = 82'b1000001100100100101100110001111100001101101101100001010100001010010111001001011000;
	ram[928] = 82'b1000001100011100000110010101100111110001110000010010100010101101110010010100000000;
	ram[929] = 82'b1000001100010011100000010100010110100011010000000101111111100111000110110111101000;
	ram[930] = 82'b1000001100001010111010101110000111011111111010110001101101000100100110110010011110;
	ram[931] = 82'b1000001100000010010101100010110111100111111011001001000010101101110001100000100001;
	ram[932] = 82'b1000001011111001110000110010100101000111001001000111001100100011111011100100010100;
	ram[933] = 82'b1000001011110001001100011101001101010111011100011000010101000101010100101011111000;
	ram[934] = 82'b1000001011101000101000100010101110100101001011011011110100101000110111111101001110;
	ram[935] = 82'b1000001011100000000101000011000110100011110100111110001001010100010100111011111000;
	ram[936] = 82'b1000001011010111100001111110010011000111000111010001111111110001110101101101001000;
	ram[937] = 82'b1000001011001110111111010100010001101001111101100000110110110110100101110100101111;
	ram[938] = 82'b1000001011000110011101000101000000011001101011001010001011110100101101111010110110;
	ram[939] = 82'b1000001010111101111011010000011100110001101100110010001101101001100010000110001000;
	ram[940] = 82'b1000001010110101011001110110100101011000110101011010101010010001100000010011100000;
	ram[941] = 82'b1000001010101100111000110111010111010010000000001101011000011010111001110101100001;
	ram[942] = 82'b1000001010100100011000010010110000010010011110000000001010101111111010111100010010;
	ram[943] = 82'b1000001010011011111000001000101110101000101101001010111110011001011001000100110001;
	ram[944] = 82'b1000001010010011011000011001010000001010011011101000000101100000110000111001110000;
	ram[945] = 82'b1000001010001010111001000100010010101101100110011111011001000010111100010111111001;
	ram[946] = 82'b1000001010000010011010001001110011101111011110111100101100000111000010001010000000;
	ram[947] = 82'b1000001001111001111011101001110001011111011111000111110111100001111100110101101111;
	ram[948] = 82'b1000001001110001011101100100001001011011011001000111100000011000010000011111100100;
	ram[949] = 82'b1000001001101000111111111000111001110011000100101001011011010011001100101101011111;
	ram[950] = 82'b1000001001100000100010101000000000011101101101010101000101101010010101001110101010;
	ram[951] = 82'b1000001001011000000101110001011010111001110101110011011011000101011110100000111000;
	ram[952] = 82'b1000001001001111101001010101000111011000000010011011000111011111011010001011101000;
	ram[953] = 82'b1000001001000111001101010011000011110000001101001000011111011011010011100111001000;
	ram[954] = 82'b1000001000111110110001101011001101100001101001000101001110010010010110000000000000;
	ram[955] = 82'b1000001000110110010110011101100010111101100110101001000001011110111111111101000000;
	ram[956] = 82'b1000001000101101111011101010000001111100101101101110100110100101111011101010100000;
	ram[957] = 82'b1000001000100101100001010000100111111111000010000100001011010111110101000100010011;
	ram[958] = 82'b1000001000011101000111010001010011010110011111010101010111010111001001111011010000;
	ram[959] = 82'b1000001000010100101101101100000001111100011011000100110111001001000010110100111101;
	ram[960] = 82'b1000001000001100010100100000110001010001101001101110100110000001100001000001000000;
	ram[961] = 82'b1000001000000011111011101111011111010000000001100001111011111010111110000100001000;
	ram[962] = 82'b1000000111111011100011011000001010100011000110111111000101001101101101110100010000;
	ram[963] = 82'b1000000111110011001011011010110000010011101100110101100110111000101110000011000011;
	ram[964] = 82'b1000000111101010110011110111001110011100010110111110111111100110010111000010111100;
	ram[965] = 82'b1000000111100010011100101101100011101001010010000010000110100000011100001011001000;
	ram[966] = 82'b1000000111011010000101111101101100101011010110111100000100100000000000100111001110;
	ram[967] = 82'b1000000111010001101111100111101000100111111010101000000100001000100111011110110011;
	ram[968] = 82'b1000000111001001011001101011010100101001000010111111100011101111110001001000000000;
	ram[969] = 82'b1000000111000001000100001000101110101010011110100011001000110001000110001111101000;
	ram[970] = 82'b1000000110111000101110111111110101011001011100111100101100010000010010111111010010;
	ram[971] = 82'b1000000110110000011010010000100110000000110101000100100100010110111110001111110101;
	ram[972] = 82'b1000000110101000000101111010111110011101000010011001000100011011001100000000000000;
	ram[973] = 82'b1000000110011111110001111110111101000011010100111001011111001101101111111011010011;
	ram[974] = 82'b1000000110010111011110011100011111110000100010110110100011010010110101001010000000;
	ram[975] = 82'b1000000110001111001011010011100100001001001100010110011101011111001010001000000000;
	ram[976] = 82'b1000000110000110111000100100001000100011001011001110110011000111000110111010000000;
	ram[977] = 82'b1000000101111110100110001110001010100011011110011001110110001011111101100000100011;
	ram[978] = 82'b1000000101110110010100010001101000100000011011100000110110011011010110001000010000;
	ram[979] = 82'b1000000101101110000010101110100000011000000001111000100010000110010010001101000101;
	ram[980] = 82'b1000000101100101110001100100101111101111111110010101010101000110000110111111111100;
	ram[981] = 82'b1000000101011101100000110100010100111111001111101100001000111011101010110011101001;
	ram[982] = 82'b1000000101010101010000011101001101101100000001011011101110001001110110100001010000;
	ram[983] = 82'b1000000101001101000000011111011000001101101101101100011111000000000101000011110011;
	ram[984] = 82'b1000000101000100110000111010110010100011011011111100100110100111010010110111000000;
	ram[985] = 82'b1000000100111100100001101111011010010100000101011100000101011010001110001111011000;
	ram[986] = 82'b1000000100110100010010111101001101011111010000101000001110001100110001101100111010;
	ram[987] = 82'b1000000100101100000100100100001010011101001101110100001111110000010000111101111000;
	ram[988] = 82'b1000000100100011110110100100001111001101111110010011100001001010001010110011011100;
	ram[989] = 82'b1000000100011011101000111101011001110001110000110011100111000011111010011010111000;
	ram[990] = 82'b1000000100010011011011101111100111110000101001100110010010010010111110010000110000;
	ram[991] = 82'b1000000100001011001110111010110111001011010110101101000111010110011101101111011011;
	ram[992] = 82'b1000000100000011000010011111000110011011001011011001100110101010101110100100000000;
	ram[993] = 82'b1000000011111010110110011100010011100001001111100001010001101001111101110100000101;
	ram[994] = 82'b1000000011110010101010110010011100000110100010111110000011100101000010011001000110;
	ram[995] = 82'b1000000011101010011111100001011110100101000000111110100101111110110100001100110101;
	ram[996] = 82'b1000000011100010010100101001011000100110000111010010101011001110010111001100100000;
	ram[997] = 82'b1000000011011010001010001010001000100100001011011101110101011010101110111010111111;
	ram[998] = 82'b1000000011010010000000000011101100001001001000101001001011110111100000001101100010;
	ram[999] = 82'b1000000011001001110110010110000001101111101110111001110010010011000000010010111111;
	ram[1000] = 82'b1000000011000001101101000001000111000010010110010110111111101000010101010011000000;
	ram[1001] = 82'b1000000010111001100100000100111010011100001001110010100111010101011011001101101001;
	ram[1002] = 82'b1000000010110001011011100001011010000000001110100011010010111000100111101001010000;
	ram[1003] = 82'b1000000010101001010011010110100011011001101000010011101111111111100000101001011000;
	ram[1004] = 82'b1000000010100001001011100100010101000100001000110000110110101110100000000000000000;
	ram[1005] = 82'b1000000010011001000100001010101100101011010001000101000000100001001011111100000001;
	ram[1006] = 82'b1000000010010000111101001001101000101011001100011111011001000001111011010000000000;
	ram[1007] = 82'b1000000010001000110110100001000110101111111001010100001001111111000000111100111000;
	ram[1008] = 82'b1000000010000000110000010001000101010101111100011010111101101011000001000110000000;
	ram[1009] = 82'b1000000001111000101010011001100010001001110000111101001110111000000111010000010001;
	ram[1010] = 82'b1000000001110000100100111010011011101000010101011111110111001111100000101010110000;
	ram[1011] = 82'b1000000001101000011111110011101111011110100001101110011111011100001001101100111000;
	ram[1012] = 82'b1000000001100000011011000101011100001001101101111110100111000001000001101100000000;
	ram[1013] = 82'b1000000001011000010110101111011111010111001110001100011101010001101001010011111001;
	ram[1014] = 82'b1000000001010000010010110001110111100100110100100000000100001011000111101010000000;
	ram[1015] = 82'b1000000001001000001111001100100010111000010111000011111000011101101000110100011111;
	ram[1016] = 82'b1000000001000000001011111111011110111111110100100001011010110101011011110010011000;
	ram[1017] = 82'b1000000000111000001001001010101010000001100000011100000111000100111000000000000000;
	ram[1018] = 82'b1000000000110000000110101110000010011011111111000001010010101010010111110100101010;
	ram[1019] = 82'b1000000000101000000100101001100101111101111001000011010100101000010110010111101011;
	ram[1020] = 82'b1000000000100000000010111101010011000110001100011111011100011100111001001101100100;
	ram[1021] = 82'b1000000000011000000001101001000111111011111111101011000111111111011010110101110111;
	ram[1022] = 82'b1000000000010000000000101101000010001110100101001010001110010000001110000000010000;
	ram[1023] = 82'b1000000000001000000000001001000000000101100000000001000000000000000000000000000000;
end
endmodule

module sqrt_load_grad_table (
    input wire [9:0] addr,
    output wire [70:0] grd,
    input wire clk,
	input wire rstn);

(* RAM_STYLE="BLOCK" *) reg [70:0] ram [1023:0];
//always @(posedge clk)
//    grd <= ram[addr];
assign grd = ram[addr];
initial begin
	ram[0] = 71'b10110100111000110000101010110110010001011011000000100010011111001011101;
	ram[1] = 71'b10110100100111110101001110100010010100101010011010111001001100110010101;
	ram[2] = 71'b10110100010110111100010101100111110010001010001111100110101000101100101;
	ram[3] = 71'b10110100000110000110001011110000000000010100010000011010100010000011000;
	ram[4] = 71'b10110011110101010010100100101000000111110100100001011001010001110100111;
	ram[5] = 71'b10110011100100100001101011111000000101100101111000100001001101100000001;
	ram[6] = 71'b10110011010011110011010101001110100111100001010000101001011111001001011;
	ram[7] = 71'b10110011000011000111100000010111110110110000111011101001001011111110101;
	ram[8] = 71'b10110010110010011110001100111111111111001011010100111111100011001101111;
	ram[9] = 71'b10110010100001110111100110101100001011011111001001111111000100100101000;
	ram[10] = 71'b10110010010001010011101101000110011111101011011110001110110100000111000;
	ram[11] = 71'b10110010000000110010001000001010000110101011100100000010110100101111001;
	ram[12] = 71'b10110001110000010011001111010011000010110001011010101000110010101110101;
	ram[13] = 71'b10110001011111110110110110010101100000100110100100111001110101000101001;
	ram[14] = 71'b10110001001111011100111100111101111100100111001001001000011011101010101;
	ram[15] = 71'b10110000111111000101100010111000110101111001100110010101110101100111001;
	ram[16] = 71'b10110000101110110000110011100110100010110010110000101111111101010111000;
	ram[17] = 71'b10110000011110011110010111001011010000000111111011100010010011100101000;
	ram[18] = 71'b10110000001110001110100100111010011111110100100110110010010010011001111;
	ram[19] = 71'b10101111111110000001010000101101000111010011000101000000100000011000000;
	ram[20] = 71'b10101111101101110110011010001111110011001010111110001110010011011010001;
	ram[21] = 71'b10101111011101101110000001001111010010101100110100011011100011111111000;
	ram[22] = 71'b10101111001101101000010001000111110111000000011010110110001111101000000;
	ram[23] = 71'b10101110111101100100110010000110101000001111100011111011111100110010001;
	ram[24] = 71'b10101110101101100011101111101000101010110010110111100101110010010011000;
	ram[25] = 71'b10101110011101100101001001011010111000011100000101000000000011110011011;
	ram[26] = 71'b10101110001101101000111111001010001101100100101000010010000111000000000;
	ram[27] = 71'b10101101111101101111011100001111100011101111010110010010000000000011000;
	ram[28] = 71'b10101101101101111000001000111111011010000001110011110011111000101000011;
	ram[29] = 71'b10101101011110000011010000110011011100110001010011111111010001000000000;
	ram[30] = 71'b10101101001110010000110011011000110010110011101101000000010111010000101;
	ram[31] = 71'b10101100111110100000100100110011100000011100110101101100111011101101001;
	ram[32] = 71'b10101100101110110010111100000011101001001000110011100011011011101111000;
	ram[33] = 71'b10101100011111000111101101001100101001001001101111101011101000000110011;
	ram[34] = 71'b10101100001111011110101100010100110011101110111011010010110001001111111;
	ram[35] = 71'b10101011111111111000000100110001110100011011110010001110001000110000011;
	ram[36] = 71'b10101011110000010011110110010001000001011001000100101001110000101111111;
	ram[37] = 71'b10101011100000110010000000011111110011010100101001100111101111000110011;
	ram[38] = 71'b10101011010001010010010111100111011010100010111111010010010101101111000;
	ram[39] = 71'b10101011000001110101000110111010111000111110110111100011011001101101001;
	ram[40] = 71'b10101010110010011010001110000111101110110011100011000100101100111000000;
	ram[41] = 71'b10101010100011000001101100111011011110110000011110100011011100111010111;
	ram[42] = 71'b10101010010011101011010111100010010100110101101011011001111001101101001;
	ram[43] = 71'b10101010000100010111011001001100101010100111111001100001000000001101011;
	ram[44] = 71'b10101001110101000101110001101000001010010001010011110000010001000001101;
	ram[45] = 71'b10101001100101110110010101000011001011100100001101011000000010111111000;
	ram[46] = 71'b10101001010110101001001110101100001010100110101011001000000011011101111;
	ram[47] = 71'b10101001000111011110011110010000111000111011100111001010111101000000000;
	ram[48] = 71'b10101000111000010101111000000001111001010101111110000001100001000000000;
	ram[49] = 71'b10101000101001001111011011101111000101100110100000100101101000011001111;
	ram[50] = 71'b10101000011010001011010100100100010011011100001101010000111101001111000;
	ram[51] = 71'b10101000001011001001100010001111011110000010010110000001111111101101101;
	ram[52] = 71'b10100111111100001001111001000100000000001011110100000011001101100001011;
	ram[53] = 71'b10100111101101001100100100001011110011110010100001010100000000001001001;
	ram[54] = 71'b10100111011110010001010111111011101111001000110000100011111111101011000;
	ram[55] = 71'b10100111001111011000011111011100011001111000111001010101101100110000011;
	ram[56] = 71'b10100111000000100001101111000100000101011111001001001101000101010000111;
	ram[57] = 71'b10100110110001101101000110100010111100111010000101011100010101000101000;
	ram[58] = 71'b10100110100010111010110000111111101100111001111111011111101110110011101;
	ram[59] = 71'b10100110010100001010100010110010101110111010100101101010101011100000111;
	ram[60] = 71'b10100110000101011100100111000001011110001101101000110010101110001110001;
	ram[61] = 71'b10100101110110110000110010000101101110100011110100000111010001011001000;
	ram[62] = 71'b10100101101000000111000011101111110101011110101111101000110111110101000;
	ram[63] = 71'b10100101011001011111100111000011010100011111011111010110010101101101000;
	ram[64] = 71'b10100101001010111010000101001001100110101001011000000000000000000000000;
	ram[65] = 71'b10100100111100010110111111101010100110000110110110111000000111100011111;
	ram[66] = 71'b10100100101101110101110100011111010010010000011111101001001010001000000;
	ram[67] = 71'b10100100011111010110111001111011001010101101001000000010110101010010001;
	ram[68] = 71'b10100100010000111010000100011100111100011011000100011000100101101011101;
	ram[69] = 71'b10100100000010011111010011110101001011011001100000100001000000000000000;
	ram[70] = 71'b10100011110100000110100111110100011101100110111110111000111001110001000;
	ram[71] = 71'b10100011100101110000001011011001010011000001010001110010101110011000000;
	ram[72] = 71'b10100011010111011011110011000101001001110001100100010010001111000100101;
	ram[73] = 71'b10100011001001001001010011011100001001101111111100000101110101101000000;
	ram[74] = 71'b10100010111010111001000010101000110011011000101101001100001100101101011;
	ram[75] = 71'b10100010101100101010110101001110101000101100011001101110000100110001001;
	ram[76] = 71'b10100010011110011110110110001001000011000001000111001110001110100010111;
	ram[77] = 71'b10100010010000010100101110110010111110010111100011000110010001010000011;
	ram[78] = 71'b10100010000010001100101010001000100001101000001010001111110110100011000;
	ram[79] = 71'b10100001110100000110110011000011001111101101010010111000010100000101001;
	ram[80] = 71'b10100001100110000010110011000010000011011010100101100111111001100001000;
	ram[81] = 71'b10100001011000000001000000000110100101010111011010001110000001011001011;
	ram[82] = 71'b10100001001010000001000011110010011001011101101100101000000011001101000;
	ram[83] = 71'b10100000111100000011010100000100100111010110101010111101010011000011001;
	ram[84] = 71'b10100000101110000111011010100001011011011011110000001000110011000111000;
	ram[85] = 71'b10100000100000001101101101000101011100111101011011101010011111101100011;
	ram[86] = 71'b10100000010010010101110101010111100000001101111000001000101010010111000;
	ram[87] = 71'b10100000000100011111111110001110001010000001000001101011010001000000000;
	ram[88] = 71'b10011111110110101100000111011010100011111010100110011001000110101011001;
	ram[89] = 71'b10011111101000111010011011110000001010101110000011110001101000011001000;
	ram[90] = 71'b10011111011011001010100100111011000000101100001011100100111011011100001;
	ram[91] = 71'b10011111001101011100100010101110001110110111011110010010001000100011000;
	ram[92] = 71'b10011110111111110000101010111101101111011111010011101001101000000001011;
	ram[93] = 71'b10011110110010000110110010011001001101000010001101110110101010100100111;
	ram[94] = 71'b10011110100100011110101101110010110101011010000000011110010100001100001;
	ram[95] = 71'b10011110010110111000100111111100010111010100001101111011110100111001000;
	ram[96] = 71'b10011110001001010100100000100111001011100010100001110100010100111101000;
	ram[97] = 71'b10011101111011110010010111100100101100110001011001001110101000100011001;
	ram[98] = 71'b10011101101110010010000001101001110000101110101101110000000011010111000;
	ram[99] = 71'b10011101100000110011101001100101101100101001010111001111100101110101000;
	ram[100] = 71'b10011101010011010111001111001010000000101111000101000100001000001110101;
	ram[101] = 71'b10011101000101111100110010001000001111000111101110110011001111101010111;
	ram[102] = 71'b10011100111000100100000111010111110100001001110111000010100111001110111;
	ram[103] = 71'b10011100101011001101100100011111001100101111010101111010001110101101111;
	ram[104] = 71'b10011100011101111000101000100011100000010110000110000100001101111000000;
	ram[105] = 71'b10011100010000100101110100000010111000101000001111101010000111000010001;
	ram[106] = 71'b10011100000011010100110000111101110111010110101101000101100110011000000;
	ram[107] = 71'b10011011110110000101011111000111111111110110111001000001111110101110101;
	ram[108] = 71'b10011011101000111000010100000001101100110111100000111000001001100011000;
	ram[109] = 71'b10011011011011101100101110111001011110001001000101110110101010001000000;
	ram[110] = 71'b10011011001110100011010000000100010111000110010010110011001011110101000;
	ram[111] = 71'b10011011000001011011100001101001001011101000111001101001011000000011000;
	ram[112] = 71'b10011010110100010101100011011011100111000011011101001011101011000000000;
	ram[113] = 71'b10011010100111010001101010110110000101010011111010100010110001100001000;
	ram[114] = 71'b10011010011010001111010111010000011001001100110101101000001100111010001;
	ram[115] = 71'b10011010001101001110111110000100011011000101101101100010010110000110111;
	ram[116] = 71'b10011010000000010000011111000100001000000111110101001100110001001000000;
	ram[117] = 71'b10011001110011010011101111010000100010110000001001100001011000010110111;
	ram[118] = 71'b10011001100110011000111001001101110101100101111110111100001001011010001;
	ram[119] = 71'b10011001011001011111110001111110010011101110101001101011001011001000001;
	ram[120] = 71'b10011001001100101000011001010101110100111010010111110001110010000000111;
	ram[121] = 71'b10011000111111110010111001110110110100111011110111111111111000101000000;
	ram[122] = 71'b10011000110010111111001000100101011111001101011001111010101010101000111;
	ram[123] = 71'b10011000100110001101010000000011000110000010010100001010011000011000001;
	ram[124] = 71'b10011000011001011101000101010101000100110000111100101110011001010010001;
	ram[125] = 71'b10011000001100101110110010111011100100011110000010110000111101000000000;
	ram[126] = 71'b10011000000000000010000011010001101100100001011010110110000011001000000;
	ram[127] = 71'b10010111110011010111010110001110001010010010100001011111111101000000000;
	ram[128] = 71'b10010111100110101110001011100010010110110000010010001001100111010010001;
	ram[129] = 71'b10010111011010000110111000010111101100101111011110001001101101011000001;
	ram[130] = 71'b10010111001101100001010001110111010101100100001000000110000110101000111;
	ram[131] = 71'b10010111000000111101010111110101011001100111001111110110010110011101011;
	ram[132] = 71'b10010110110100011011010100101110000011011000001001010011001101110011000;
	ram[133] = 71'b10010110100111111010111101101100010010001111001100101000001100000111111;
	ram[134] = 71'b10010110011011011100010010100100010011000100000001011100010100100111000;
	ram[135] = 71'b10010110001110111111010011001010010100001001011111111111111011001111011;
	ram[136] = 71'b10010110000010100100001001111000001111110111111000000001011001100011111;
	ram[137] = 71'b10010101110110001010101011111011100010000010000111000101101001011100001;
	ram[138] = 71'b10010101101001110010111001001000011101011000001101110010110111101111001;
	ram[139] = 71'b10010101011101011100110001010011010110000100111110101011101111111100111;
	ram[140] = 71'b10010101010001001000010100010000100001101101110110110101100111110110011;
	ram[141] = 71'b10010101000100110101101100010111000111111001010001010000011011101011000;
	ram[142] = 71'b10010100111000100100101110110111100110011000011100011011110010000010111;
	ram[143] = 71'b10010100101100010101010001000100110000100100000000011011001111001110101;
	ram[144] = 71'b10010100100000000111100111110110110100000000010010010010010000010101000;
	ram[145] = 71'b10010100010011111011101000100000000001111101000001010011101110000010101;
	ram[146] = 71'b10010100000111110001010010110100111000101001001011011011100000011011000;
	ram[147] = 71'b10010011111011101000100110101001110111101101100100100101100010011111101;
	ram[148] = 71'b10010011101111100001101110010010001110111110111001110001111111000110011;
	ram[149] = 71'b10010011100011011100010100100100011110101111101111101111001111110011000;
	ram[150] = 71'b10010011010111011000100011110100011110010001001001010101101100110110111;
	ram[151] = 71'b10010011001011010110011011110110110010110010001001000110000110011111000;
	ram[152] = 71'b10010010111111010110000110111100011111110000011110011010001000111000000;
	ram[153] = 71'b10010010110011010111010000000000101111001101010110101110110110011111111;
	ram[154] = 71'b10010010100111011010000001010101001011110010000101011010101101000000000;
	ram[155] = 71'b10010010011011011110100101001001010000010011101011011011110011000000000;
	ram[156] = 71'b10010010001111100100100110011011100100110001101101001010001000010010101;
	ram[157] = 71'b10010010000011101100001111011100001011000000001100110011101001000000000;
	ram[158] = 71'b10010001110111110101011111111111110001111100101110000000110010101011001;
	ram[159] = 71'b10010001101100000000010111111011001001111101010011000101101000000000000;
	ram[160] = 71'b10010001100000001100110111000011000100110000010101110011111010001000101;
	ram[161] = 71'b10010001010100011010111101001100010101011100100000001101111000000000000;
	ram[162] = 71'b10010001001000101010101010001011110000100000100101011001100011100011001;
	ram[163] = 71'b10010000111100111011110011011111111011010000000101000101101100100110111;
	ram[164] = 71'b10010000110001001110101101101010110001101010100000110111111111011000000;
	ram[165] = 71'b10010000100101100011000011110101001110110010100011100110000001000011000;
	ram[166] = 71'b10010000011001111001000000001010011100111110000011011101000100101011000;
	ram[167] = 71'b10010000001110010000100010011111010111010111000111100101110000111000000;
	ram[168] = 71'b10010000000010101001101010101000111010011111010110001001110011000000000;
	ram[169] = 71'b10001111110111000100011000011100000100001111101101001011010111110101000;
	ram[170] = 71'b10001111101011100000100001011011011011101101010100000110011101100100001;
	ram[171] = 71'b10001111011111111110001111101111100000001001101111111001010111100111000;
	ram[172] = 71'b10001111010100011101100011001101010011010111110001001010010001110000001;
	ram[173] = 71'b10001111001000111110011011101001111000100001000100110111110101010101000;
	ram[174] = 71'b10001110111101100000101110101010001000100011011010101001000111000000000;
	ram[175] = 71'b10001110110010000100100110010100011010111001110101111100111100111000000;
	ram[176] = 71'b10001110100110101010000010011101110110100110100110110011101010011011000;
	ram[177] = 71'b10001110011011010000111000101101000001010110110011000001110010010001101;
	ram[178] = 71'b10001110001111111001011101010100101101000110000100111001000101001010011;
	ram[179] = 71'b10001110000100100011011011101101100010010000011101101110101100001011000;
	ram[180] = 71'b10001101111001001110110011101110010101011011010101101011001101101011000;
	ram[181] = 71'b10001101101101111011101111011010010011110111110101010000110110011000000;
	ram[182] = 71'b10001101100010101010001110100110101100010110100010011010101111000000000;
	ram[183] = 71'b10001101010111011010010001001000101110111101111011110000101110011101000;
	ram[184] = 71'b10001101001100001011101100101010111101000111011100111000010111101100001;
	ram[185] = 71'b10001101000000111110100001000100010000110111111011111101110001001100101;
	ram[186] = 71'b10001100110101110011000010011110111011110000100011001111000000000000000;
	ram[187] = 71'b10001100101010101000111100011100011010000101111101001101011001000000000;
	ram[188] = 71'b10001100011111100000001110110011101001010000110100100010001100100001101;
	ram[189] = 71'b10001100010100011001000011100011101100000101000110100011011101000000000;
	ram[190] = 71'b10001100001001010011011010100001111011011101000010001111001001011100001;
	ram[191] = 71'b10001011111110001111001001011100110001011011011101100100110011001011111;
	ram[192] = 71'b10001011110011001100010000001011001111101011100011011111100111110001000;
	ram[193] = 71'b10001011101000001011000010110000010001001100110000010010101110011000000;
	ram[194] = 71'b10001011011101001011000010101111011111010110000000101101101110000101000;
	ram[195] = 71'b10001011010010001100100100001011010101011011010011001011011110110111000;
	ram[196] = 71'b10001011000111001111100110111001010011110001010111011010000101000000000;
	ram[197] = 71'b10001010111100010100000000101011000111001110100010011110001000111010111;
	ram[198] = 71'b10001010110001011001111011011011001010111100100111011111000110011000000;
	ram[199] = 71'b10001010100110100001001100111100010001100101101100100010000001010011000;
	ram[200] = 71'b10001010011011101001110101000101100101010101110101010010000100011111101;
	ram[201] = 71'b10001010010000110011111101101111111111101010110100110011001101000101000;
	ram[202] = 71'b10001010000101111111011100101111111011011100010001110011100100101000000;
	ram[203] = 71'b10001001111011001100011011111101010001010100100000101100110110101000000;
	ram[204] = 71'b10001001110000011010110001001101100001011011000000111010001010000101001;
	ram[205] = 71'b10001001100101101010100110010111100011110100011011011000101110001000000;
	ram[206] = 71'b10001001011010111011110001010001111101101001100111111110111111101000000;
	ram[207] = 71'b10001001010000001110010001110100000000011010000011000110011001101111001;
	ram[208] = 71'b10001001000101100010000111110100111110100011010111000111000100101011011;
	ram[209] = 71'b10001000111010110111011101001001101111011100110111010001010111011111011;
	ram[210] = 71'b10001000110000001110000111101011000001011101011100111000010001000000000;
	ram[211] = 71'b10001000100101100110010001001100101011111111000011100110011100011101011;
	ram[212] = 71'b10001000011010111111101111101000100001101111100110000011100011100111011;
	ram[213] = 71'b10001000010000011010100010110101111010010110010011011011110011000000000;
	ram[214] = 71'b10001000000101110110101010101100001110011000001011001100101010111001000;
	ram[215] = 71'b10000111111011010100010000111101010101110010010000101001100100111001000;
	ram[216] = 71'b10000111110000110011001011100101001011001100000100001100100000101000111;
	ram[217] = 71'b10000111100110010011011010011011001010001101001010101001001111100100001;
	ram[218] = 71'b10000111011011110101000111001111101011110010010101011000010001101010001;
	ram[219] = 71'b10000111010001011000001000000000001111111100010010110010110011011011000;
	ram[220] = 71'b10000111000110111100010010101100011010000010111100100111010111011011111;
	ram[221] = 71'b10000110111100100010000100110011011011100001100100100011011100000111111;
	ram[222] = 71'b10000110110010001001000000100101000011000111010111000010000011010111011;
	ram[223] = 71'b10000110100111110001001111110000101101100110101111001011011011011000000;
	ram[224] = 71'b10000110011101011010111100000011110111001010000100000100111001001000011;
	ram[225] = 71'b10000110010011000101111011011111001000111101100011100010001101101001111;
	ram[226] = 71'b10000110001000110010001101111010000111100010100100011101101101000000000;
	ram[227] = 71'b10000101111110011111110011001100011000010111001111011001110001101011000;
	ram[228] = 71'b10000101110100001110110101000001011010110011011001010110101110101101000;
	ram[229] = 71'b10000101101001111110111111101000100100010000100101010001110101101001000;
	ram[230] = 71'b10000101011111110000100110100000101110111111110001111000000000000000000;
	ram[231] = 71'b10000101010101100011010101111011010010100010010111111010001101011001000;
	ram[232] = 71'b10000101001011010111100001010101001011000000010010100110110010001101000;
	ram[233] = 71'b10000101000001001100111110110011001010110011100111011001101101010010111;
	ram[234] = 71'b10000100110111000011101110001100111110001011100000000110001100000111001;
	ram[235] = 71'b10000100101100111011101111011010010010010011010010101011001000000000000;
	ram[236] = 71'b10000100100010110101000010010010110101010010011100101110111111111000000;
	ram[237] = 71'b10000100011000101111100110101110010110001100011110111100000111110110101;
	ram[238] = 71'b10000100001110101011011100100100100101000000111000011101001110110111011;
	ram[239] = 71'b10000100000100101000100011101101010010101011000010011010011010001111000;
	ram[240] = 71'b10000011111010100110111100000000010001000010001011010110010111001111000;
	ram[241] = 71'b10000011110000100110101111000010101111000010101101111000011001001000000;
	ram[242] = 71'b10000011100110100111101001010001001000101110100101111011110010100111000;
	ram[243] = 71'b10000011011100101001110100010001001110010110100111000101100100101100101;
	ram[244] = 71'b10000011010010101101001111111010110101100000101000000010111111100110001;
	ram[245] = 71'b10000011001000110001111100000101110100101101111110010011011101101101000;
	ram[246] = 71'b10000010111110110111111000101010000011011011011001100111111001000000000;
	ram[247] = 71'b10000010110100111111000101011111011010000000111111100010010110011010011;
	ram[248] = 71'b10000010101011000111100010011101110001110010000110110110000111001001011;
	ram[249] = 71'b10000010100001010001001111011101000100111101010011001000000000000000000;
	ram[250] = 71'b10000010010111011100001100010101001110101100010000001111000110101001000;
	ram[251] = 71'b10000010001101101000011000111110001011000011101101110101110100110111001;
	ram[252] = 71'b10000010000011110101110101001111110111000011011010111011010001110011101;
	ram[253] = 71'b10000001111010000100010111011010101010000010010010101101000000011011101;
	ram[254] = 71'b10000001110000010100001000111111000111000001111100110111000001001101000;
	ram[255] = 71'b10000001100110100101010011011011110110100111010000100011100101100001101;
	ram[256] = 71'b10000001011100110111100011011011001000101001100111111010001100001000000;
	ram[257] = 71'b10000001010011001011000010011100000110010100100100001100110011000000000;
	ram[258] = 71'b10000001001001011111110000010110110001111110111000111110000101110010001;
	ram[259] = 71'b10000000111111110101100011011110100000100001101011000000100101010111000;
	ram[260] = 71'b10000000110110001100101110110101010001011010110001010001101001011010001;
	ram[261] = 71'b10000000101100100100111111001010001011011011101010010110000011000000000;
	ram[262] = 71'b10000000100010111110011101111010000010110011101010001001011010001000000;
	ram[263] = 71'b10000000011001011001001010111100111110010100000100110110110000000001101;
	ram[264] = 71'b10000000001111110101000110001011000101101000011010000011100000100010011;
	ram[265] = 71'b10000000000110010010000101111010101001011011101001100101111000001011101;
	ram[266] = 71'b01111111111100110000011101001000000001010010000001000100100000001011101;
	ram[267] = 71'b01111111110011001111111000101000000101111001100001010101000001110111001;
	ram[268] = 71'b01111111101001110000011000010100011101000010100000111111101101000010001;
	ram[269] = 71'b01111111100000010010001111000110101011100000011011101101111111100111111;
	ram[270] = 71'b01111111010110110101001001110110100001101000111110000010110101001110001;
	ram[271] = 71'b01111111001101011001010001111100101010011110110010100111100101000000000;
	ram[272] = 71'b01111111000011111110100111010001010100101001110001010100000000001000000;
	ram[273] = 71'b01111110111010100101000000001110101000011010110010101111011011001000000;
	ram[274] = 71'b01111110110001001100100110001011111001001100110101111000010111110011001;
	ram[275] = 71'b01111110100111110101011001000001011000001011000100000111100010011101011;
	ram[276] = 71'b01111110011110011111001111001010101001101000011111110011000110111100001;
	ram[277] = 71'b01111110010101001010010001111101101001110010010110101000110001101000000;
	ram[278] = 71'b01111110001011110110100001010010101100010110011111111011011011011000000;
	ram[279] = 71'b01111110000010100011110011100110110001001111001101011100111001000000000;
	ram[280] = 71'b01111101111001010010010010001110011101110101110001110010100111101011001;
	ram[281] = 71'b01111101110000000001111101000010001000011010001110101010110101001101111;
	ram[282] = 71'b01111101100110110010101010100000001100000011001111011111010001100001001;
	ram[283] = 71'b01111101011101100100100011111011110111101111111101100101010101000000000;
	ram[284] = 71'b01111101010100010111101001001101100100010010000001101111100001111000000;
	ram[285] = 71'b01111101001011001011110000110101000111100001101111101010010111101000000;
	ram[286] = 71'b01111101000010000001000100000100011010011101110101000011110110101010001;
	ram[287] = 71'b01111100111000110111011001011100001111001110000101101001111001111001000;
	ram[288] = 71'b01111100101111101110111010001101100101100110110011111011010111000000000;
	ram[289] = 71'b01111100100110100111011100111010001011110011110010001001100111110001000;
	ram[290] = 71'b01111100011101100001001010110010001000101001111100100110100001000110001;
	ram[291] = 71'b01111100010100011100000011101101111010101011110010111111110110011111101;
	ram[292] = 71'b01111100001011010111111110010000101001111001100000100101000000111100101;
	ram[293] = 71'b01111100000010010100111010010100001101101001001001111000010101000101001;
	ram[294] = 71'b01111011111001010011000001000110111011010010100110110101111001100101000;
	ram[295] = 71'b01111011110000010010010010100001010100100111001111000000000000000000000;
	ram[296] = 71'b01111011100111010010100101001000011000101001110010011011110001111101000;
	ram[297] = 71'b01111011011110010100000010001001001000001101100110100000010111010001001;
	ram[298] = 71'b01111011010101010110100000001001011101100101010100011010111110011000000;
	ram[299] = 71'b01111011001100011001111111000011010100001001110011001101010011101011011;
	ram[300] = 71'b01111011000011011110101000000010011000011010001010110000001001100011111;
	ram[301] = 71'b01111010111010100100011010111111010000111100011000000000000000000000000;
	ram[302] = 71'b01111010110001101011001110100001101110000001000110001100000010001011101;
	ram[303] = 71'b01111010101000110011000010100011101101101100101101111100000110110111000;
	ram[304] = 71'b01111010011111111100000000001111001100101111001111000000110111111000000;
	ram[305] = 71'b01111010010111000101111110001101010011010101111010111000111111000111000;
	ram[306] = 71'b01111010001110010001000101100111000110101001011000001111001001010011101;
	ram[307] = 71'b01111010000101011101001101000110101001010100000010101001000000000000000;
	ram[308] = 71'b01111001111100101010010100100101111100101011110000111111000001110011111;
	ram[309] = 71'b01111001110011111000100101001100110010101110001000001001111010011111011;
	ram[310] = 71'b01111001101011000111111110110011111001000111100111000101110100011000000;
	ram[311] = 71'b01111001100010011000001110111010001111011011011110011000010111000000000;
	ram[312] = 71'b01111001011001101001100111110100000100110110000001110100010101111011001;
	ram[313] = 71'b01111001010000111100001001011010001001010111010001001011001111110011111;
	ram[314] = 71'b01111001001000001111100001001110000111110001111100011100000111000000000;
	ram[315] = 71'b01111000111111100100000001100001101000001001001010111101101101110011000;
	ram[316] = 71'b01111000110110111001101010001101011100101111111110100100000101000101001;
	ram[317] = 71'b01111000101110010000001000110101111010110111110110100001100101000011111;
	ram[318] = 71'b01111000100101100111101111101010000100001010100101100100100111011101000;
	ram[319] = 71'b01111000011101000000011110100010101101001101110000110111100011000101000;
	ram[320] = 71'b01111000010100011010000011000110110101000000111110110010000000111110101;
	ram[321] = 71'b01111000001011110100101111100010110111100100011101100001101111011011101;
	ram[322] = 71'b01111000000011010000100011101111101011101111110111000001110100110001000;
	ram[323] = 71'b01110111111010101101001101010110111001100000011000010111011010110001000;
	ram[324] = 71'b01110111110010001010111110100010010111111100010011101101000000110110111;
	ram[325] = 71'b01110111101001101001101110000100001111101011011000001101011000000000000;
	ram[326] = 71'b01110111100001001001011011110110101101100010101010100110101011010100101;
	ram[327] = 71'b01110111011000101010010000111001111000010001111011110000101100011101111;
	ram[328] = 71'b01110111010000001100000100000001001101100000011101111110100111010011101;
	ram[329] = 71'b01110111000111101110110101000110111011111100011011000111001101001111111;
	ram[330] = 71'b01110110111111010010100100000101010010111001101110011111001100011000101;
	ram[331] = 71'b01110110110110110111010000110110100010010010000010010001101000100111111;
	ram[332] = 71'b01110110101110011101000100011000101010101000001000000000010111101011000;
	ram[333] = 71'b01110110100110000011110101100001010110010010101001101001011101100110001;
	ram[334] = 71'b01110110011101101011100100001010110111000011101011101000000000000000000;
	ram[335] = 71'b01110110010101010100010000001111011111010010110110001111011001011101011;
	ram[336] = 71'b01110110001100111110000010101011100100111011001010111011010010100010011;
	ram[337] = 71'b01110110000100101000101001010100111010011000001111001011111011101011000;
	ram[338] = 71'b01110101111100010100010110001001011110100111111110101000011111001011000;
	ram[339] = 71'b01110101110100000001000000000001100011100001011010100110000000001101000;
	ram[340] = 71'b01110101101011101110100110110111011110011110110010100111100111001001000;
	ram[341] = 71'b01110101100011011101001010100101100101011111101010000010001011111111000;
	ram[342] = 71'b01110101011011001100101011000110001111001000110101010110110000110111000;
	ram[343] = 71'b01110101010010111101010001010010111000001010010101111000110000011111011;
	ram[344] = 71'b01110101001010101110110100000101111100111010110101011000001111111000000;
	ram[345] = 71'b01110101000010100001001010011011100101111111110011011011010011000000000;
	ram[346] = 71'b01110100111010010100100110001011000110111010110101101011000010011101001;
	ram[347] = 71'b01110100110010001000111110010000001110100100111110101100110000101111000;
	ram[348] = 71'b01110100101001111110010010100101010111001001001011100011100101111010111;
	ram[349] = 71'b01110100100001110100100011000100111011010111010111111011110100101000000;
	ram[350] = 71'b01110100011001101011101111101001010110100100011011100110110001010011101;
	ram[351] = 71'b01110100010001100011111000001101000100101010000111110110110100110101000;
	ram[352] = 71'b01110100001001011100111100101010100010000111000100111011101010010001011;
	ram[353] = 71'b01110100000001010111000101110111000110011000100011010010100001101110001;
	ram[354] = 71'b01110011111001010010000001110110111111110010100111100111001100111001000;
	ram[355] = 71'b01110011110001001101111001100000000001011111000010000011111010011000111;
	ram[356] = 71'b01110011101001001010110101100110010101001111011100100000110001000100001;
	ram[357] = 71'b01110011100001001000100100010000101010000000111111001011101010100111000;
	ram[358] = 71'b01110011011001000111010111001100011011011010101101000000000000000000000;
	ram[359] = 71'b01110011010001000110111100100010000011000110110110001001011100000101101;
	ram[360] = 71'b01110011001001000111100101111101010100011011011000111110010111000001111;
	ram[361] = 71'b01110011000001001001000001101000010011011100000100001010000001011000000;
	ram[362] = 71'b01110010111001001011011000010101111110010010011110001010101000000110101;
	ram[363] = 71'b01110010110001001110110010110111101010110100000011001010110111001001011;
	ram[364] = 71'b01110010101001010010111111011001111100000110011011100010000101111000000;
	ram[365] = 71'b01110010100001011000001111100100100010001000111000111100101111001101000;
	ram[366] = 71'b01110010011001011110010001100101101001101001100011100010000111101100011;
	ram[367] = 71'b01110010010001100101001110001110010000100111011010110101101000000000000;
	ram[368] = 71'b01110010001001101101000101011000111100101001011011111000000001111011001;
	ram[369] = 71'b01110010000001110101110111000000010011111010101111100010000000111011000;
	ram[370] = 71'b01110001111001111111100010111110111101001010101000000011100010011010111;
	ram[371] = 71'b01110001110010001010001001001111011111101100011110100011011001011000000;
	ram[372] = 71'b01110001101010010101101001101100100011010111110000011110111101000101101;
	ram[373] = 71'b01110001100010100010000100010000110000100111111101001010000011010001000;
	ram[374] = 71'b01110001011010101111011000110110110000011100100011001111000101010101011;
	ram[375] = 71'b01110001010010111101011110100111010000010111010010101101111111111010111;
	ram[376] = 71'b01110001001011001100100111000001001100001110000111110011000000000000000;
	ram[377] = 71'b01110001000011011100100000011011110000001111110010010000101101111000000;
	ram[378] = 71'b01110000111011101101010011100011100011100101110100010011100010111000000;
	ram[379] = 71'b01110000110011111111000000010011010001111011111000000000000000000000000;
	ram[380] = 71'b01110000101100010001100110100101100111100001011000010101000101000000000;
	ram[381] = 71'b01110000100100100101000110010101010001001001011110101101100001101000000;
	ram[382] = 71'b01110000011100111001011111011100111100001011000000100001010010001000000;
	ram[383] = 71'b01110000010101001110101001001000100110111001001100111010101010101100111;
	ram[384] = 71'b01110000001101100100110100110000111000011001001011111011100111100001111;
	ram[385] = 71'b01110000000101111011110000110011011001110010010111000001010111101101000;
	ram[386] = 71'b01101111111110010011100101111001101010001010000000110011001101010111001;
	ram[387] = 71'b01101111110110101100001011010001001111010000001000000010000011000010011;
	ram[388] = 71'b01101111101111000101110010001111100111011100010011101111000111001001000;
	ram[389] = 71'b01101111100111100000001001010101101000011111000001101001100001111000000;
	ram[390] = 71'b01101111011111111011011001001011001110001110100010011100111010011101000;
	ram[391] = 71'b01101111011000010111100001101011001010110010111001010101001100111000000;
	ram[392] = 71'b01101111010000110100100010110000010000110111011101110010010000101001000;
	ram[393] = 71'b01101111001001010010010011101010100000010101001101000101000111000110011;
	ram[394] = 71'b01101111000001110001000101101010101100101011000011101010110010000111001;
	ram[395] = 71'b01101110111010010000100111010110011100100000001000100010000001011101000;
	ram[396] = 71'b01101110110010110000111000101001101111100100111000101000101101100111000;
	ram[397] = 71'b01101110101011010010001010110011000100110101011011111100000001000000111;
	ram[398] = 71'b01101110100011110100001100011010011010010011001001100000101101101011011;
	ram[399] = 71'b01101110011100010111000110000100001110100111110010100000100111101101011;
	ram[400] = 71'b01101110010100111010110111101011011000101001110000011100111010110110111;
	ram[401] = 71'b01101110001101011111011000100011000011101101111000001111011110001111000;
	ram[402] = 71'b01101110000110000100110001001110100101010100111001110000010000010001001;
	ram[403] = 71'b01101101111110101011000001101000110101110111000001101011100011000000000;
	ram[404] = 71'b01101101110111010010001001101100101110001111010101010001010110111100011;
	ram[405] = 71'b01101101101111111010000000101110111110101010000111101111100110000100001;
	ram[406] = 71'b01101101101000100010101111010001011011100111101101001000101100100010011;
	ram[407] = 71'b01101101100001001100001100101001100111011111011011100110111111000000000;
	ram[408] = 71'b01101101011001110110101001111101100101111101010001101000011111011101000;
	ram[409] = 71'b01101101010010100001101101011001010011110101101000001110001011101111000;
	ram[410] = 71'b01101101001011001101110000100110101011101100100011100011100000000100111;
	ram[411] = 71'b01101101000011111010100010010111110100011001001101001111000101010001011;
	ram[412] = 71'b01101100111100101000001011001100010001111000111010110011101101010101011;
	ram[413] = 71'b01101100110101010110101010111111000001101010000011000000000011110000111;
	ram[414] = 71'b01101100101110000101111001001000010100101110001100100110011110111111000;
	ram[415] = 71'b01101100100110110101110101100100010010100011010000001111000101000000000;
	ram[416] = 71'b01101100011111100110110001010010111011101111111001011100011100101000111;
	ram[417] = 71'b01101100011000011000011011001010111110101011101101010010000110000011001;
	ram[418] = 71'b01101100010001001010111011101001101111111110101100101110101110010111111;
	ram[419] = 71'b01101100001001111110001010001001011100010101000110111111000111000000000;
	ram[420] = 71'b01101100000010110010001111000110101000110100001100110011010100010001101;
	ram[421] = 71'b01101011111011100111000001111100010011010101100001000100000010000001101;
	ram[422] = 71'b01101011110100011100101011000110010001100011110110100001001110101101001;
	ram[423] = 71'b01101011101101010011000010000000010010011101100011011000000000000000000;
	ram[424] = 71'b01101011100110001010010111100100010111110110101100001101100001011000000;
	ram[425] = 71'b01101011011111000010010010010000110010110100011100110100011000110101000;
	ram[426] = 71'b01101011010111111011001011011101011001100010111111010010100101010110101;
	ram[427] = 71'b01101011010000110100101001101010101101110011100111101101000010000001000;
	ram[428] = 71'b01101011001001101111000110001110010111000000110110101100101110111000000;
	ram[429] = 71'b01101011000010101010010000001000001011001000011111010011010001101101001;
	ram[430] = 71'b01101010111011100110000111010100010111011111101111001010011000101001001;
	ram[431] = 71'b01101010110100100010110100001011011110000101010111000110100010001100101;
	ram[432] = 71'b01101010101101100000010110101000100101101010010110001100101110111011101;
	ram[433] = 71'b01101010100110011110100110001011010000101001101101001110101000000000000;
	ram[434] = 71'b01101010011111011101100010101111101101111001011111101101010000111111000;
	ram[435] = 71'b01101010011000011101010100101101000010000111101111000011011000000000000;
	ram[436] = 71'b01101010010001011101111011111110010101111110111110000100011111101011000;
	ram[437] = 71'b01101010001010011111010000000100101100010100100010000100010010011011111;
	ram[438] = 71'b01101010000011100001010000111100010101011110111010001011010011110100011;
	ram[439] = 71'b01101001111100100100000110111010111001011100001000110000110010111100011;
	ram[440] = 71'b01101001110101100111110001111011100010101111110101010000000110110011111;
	ram[441] = 71'b01101001101110101100000001001000001011110001010011101001111101101011101;
	ram[442] = 71'b01101001100111110001001101100110111111011011010010111100111000000000000;
	ram[443] = 71'b01101001100000110111000110100010010000011000010010000000010101011111000;
	ram[444] = 71'b01101001011001111101101011110110010001001110101000011100010100000101111;
	ram[445] = 71'b01101001010011000101000101110110011111110001011000100001110101001000000;
	ram[446] = 71'b01101001001100001101001100000111010101110011101001011000000001111000000;
	ram[447] = 71'b01101001000101010110000110111011100011010100111010011000101011000000000;
	ram[448] = 71'b01101000111110011111101101111000010001100011011011101110101001010100111;
	ram[449] = 71'b01101000110111101010000000111001110100111010000010010100010011011001001;
	ram[450] = 71'b01101000110000110101001000010001111000110110110011101010101111010111111;
	ram[451] = 71'b01101000101010000000111011100110101101011110011101111001011101000000000;
	ram[452] = 71'b01101000100011001101100011001001010000101111011000100100110010000101101;
	ram[453] = 71'b01101000011100011010110110100000100001110101000100011010111000101111101;
	ram[454] = 71'b01101000010101101000110101101000110110111110001100111000111111000000000;
	ram[455] = 71'b01101000001110110111101000110010001010000101011100001010001011111001111;
	ram[456] = 71'b01101000001000000111001111110111101101000111000110000011110011001101000;
	ram[457] = 71'b01101000000001010111011010001111000111100111011111110001110111111110111;
	ram[458] = 71'b01100111111010101000011000011010110011000111000011000010100101000000000;
	ram[459] = 71'b01100111110011111010001010010110000010110111101111011000010110000110101;
	ram[460] = 71'b01100111101101001100011111011000101001000111100101101000111100101000000;
	ram[461] = 71'b01100111100110011111101000000010110111000000110110101111110000011111111;
	ram[462] = 71'b01100111011111110011100100010000000001001010111101111100111001010111000;
	ram[463] = 71'b01100111011001001000001011101010110000010011111101011001000000000000000;
	ram[464] = 71'b01100111010010011101011110001111011110010000011010001010101000110001101;
	ram[465] = 71'b01100111001011110011011011111010100101001001100101011100000010001010101;
	ram[466] = 71'b01100111000101001010001100111000000111110000100000010111010011111111001;
	ram[467] = 71'b01100110111110100001101000110100001011010010001011101000010001000000000;
	ram[468] = 71'b01100110110111111001101111101011001010111011001111010000011011101101000;
	ram[469] = 71'b01100110110001010010101001101000000110101010110000010100101000000000000;
	ram[470] = 71'b01100110101010101100001110011000001000110001111001001010111001110101001;
	ram[471] = 71'b01100110100100000110011101110111101101100000011011011000111001111011101;
	ram[472] = 71'b01100110011101100001100000010000110010010100110100010011001110111101101;
	ram[473] = 71'b01100110010110111101001101010001100110010010100111010100110001000000000;
	ram[474] = 71'b01100110010000011001100100110110100110101100100010010110100110011111000;
	ram[475] = 71'b01100110001001110110100110111100010001001001110001100110101001000100111;
	ram[476] = 71'b01100110000011010100011011101011001010110101111011101110000010101000000;
	ram[477] = 71'b01100101111100110010111010110010111110000101001110000101100000101000000;
	ram[478] = 71'b01100101110110010010000100010000001001100001011111111101101001101100111;
	ram[479] = 71'b01100101101111110010000000001010010000011101100101000001010111111111000;
	ram[480] = 71'b01100101101001010010100110010010000001010111001110000101111001000000000;
	ram[481] = 71'b01100101100010110011110110100011111011111010110000010011110011110101101;
	ram[482] = 71'b01100101011100010101110000111100100000001000110101101000101110100011101;
	ram[483] = 71'b01100101010101111000010101011000001110010110011011100110110111000000000;
	ram[484] = 71'b01100101001111011011101011111100111100100011111100011101000101010101111;
	ram[485] = 71'b01100101001000111111101100011101001010001010001000000111001100001111001;
	ram[486] = 71'b01100101000010100100010110110101011000100000000100110101101111111011000;
	ram[487] = 71'b01100100111100001001101011000010001001010001000111000111111010001011000;
	ram[488] = 71'b01100100110101101111110001000111111011100100101100000111001101111101000;
	ram[489] = 71'b01100100101111010110011000110011000001011111001011001000111000000000000;
	ram[490] = 71'b01100100101000111101110010001111100001111100110011101010011010110101000;
	ram[491] = 71'b01100100100010100101110101010010000010110110111111001001001101000010111;
	ram[492] = 71'b01100100011100001110101001111101101100111001100100010100100111000000000;
	ram[493] = 71'b01100100010101111000000000000001100011001001010101011001100011110010011;
	ram[494] = 71'b01100100001111100010000111100110111110011100101111101011010011110001000;
	ram[495] = 71'b01100100001001001100111000100011111101110100011000101110011010111000000;
	ram[496] = 71'b01100100000010111000010010110101000101111011010010011010101110110001001;
	ram[497] = 71'b01100011111100100100010110010110111011110000011111110000001000000001001;
	ram[498] = 71'b01100011110110010001000011000110000100100111000011100111010110111000000;
	ram[499] = 71'b01100011101111111110100001000011010010111100110101100011001111101111011;
	ram[500] = 71'b01100011101001101100100000000010011101010011111101011100011010011000000;
	ram[501] = 71'b01100011100011011011010000001000001110000001110100010011011000001101001;
	ram[502] = 71'b01100011011101001010101001001100111110110111101011100111000111100011001;
	ram[503] = 71'b01100011010110111010101011001101010110110001100100010000000000111000000;
	ram[504] = 71'b01100011010000101011010110000101111100111111010111010000110110101001000;
	ram[505] = 71'b01100011001010011100101001110011011001000100110100101000001100110110011;
	ram[506] = 71'b01100011000100001110100110010010010010111001100010000001110101010110111;
	ram[507] = 71'b01100010111110000001010011100000110010111011000000001001000101110010111;
	ram[508] = 71'b01100010110111110100100001011000001011100111100010001000001000111111001;
	ram[509] = 71'b01100010110001101000011111110111110000111101100010101110101000100101111;
	ram[510] = 71'b01100010101011011101000110111010101011110110111011000100100111000000000;
	ram[511] = 71'b01100010100101010010001110011101011011001000010110010110100111100111011;
	ram[512] = 71'b01100010011111001000000110011101010011010000101011011011010101011001000;
	ram[513] = 71'b01100010011000111110100110110110011110010100111110010011100010001000000;
	ram[514] = 71'b01100010010010110101101111100101100110110000000100011011111001000101001;
	ram[515] = 71'b01100010001100101101101000100110001100110000110100010000000000001001000;
	ram[516] = 71'b01100010000110100110000001110110111011001010010100101110111011100110101;
	ram[517] = 71'b01100010000000011111000011010011101000000010110001011111100111100010011;
	ram[518] = 71'b01100001111010011000101100111000111111000011100010001010010100011000000;
	ram[519] = 71'b01100001110100010011000110100001001100111011011101110010011111010010001;
	ram[520] = 71'b01100001101110001110000000001101100111001111111001100111011111000000000;
	ram[521] = 71'b01100001101000001001100001111000110000011111111011011111000100100001000;
	ram[522] = 71'b01100001100010000101110011011011110111000100100010100011001000000000000;
	ram[523] = 71'b01100001011100000010100100111010010000000011111000011011000000000000000;
	ram[524] = 71'b01100001010110000000000110001001010111000001000010000011110010101000000;
	ram[525] = 71'b01100001001111111110000111001101110101110000111111100101110001111101000;
	ram[526] = 71'b01100001001001111100110111111011110100011100110010100001110101001000000;
	ram[527] = 71'b01100001000011111100001000011001010001011010010111111000000000000000000;
	ram[528] = 71'b01100000111101111100001000011001000001100110011101000101000000000000000;
	ram[529] = 71'b01100000110111111100101000000010010111101010000011101010001101000001000;
	ram[530] = 71'b01100000110001111101110111000110110101100011010011000110110101000000000;
	ram[531] = 71'b01100000101011111111100101101111000010000000011010011001101000000000000;
	ram[532] = 71'b01100000100110000010000011101011001100001110100111111001101101111000000;
	ram[533] = 71'b01100000100000000101000001000101001110110011100010010001101010101101000;
	ram[534] = 71'b01100000011010001000101101101100000110011001001010010100110010111000000;
	ram[535] = 71'b01100000010100001100111001101011000001001110101001111010001000000000000;
	ram[536] = 71'b01100000001110010001110100101111101001101000011110100100100001000000000;
	ram[537] = 71'b01100000001000010111001111000110100001010001100010001010001010000001000;
	ram[538] = 71'b01100000000010011101010000100100101100000101110010011001010000011111111;
	ram[539] = 71'b01011111111100100011111001000110111100000101111101101000111110011111111;
	ram[540] = 71'b01011111110110101011010000100000101110101010111011000110010000100011011;
	ram[541] = 71'b01011111110000110011000111000001001011101110100111000101100011111011001;
	ram[542] = 71'b01011111101010111011100100011100000101110101001011101111001101011001000;
	ram[543] = 71'b01011111100101000100101000101110010000001100000001100111001110101111000;
	ram[544] = 71'b01011111011111001110010011110100011110010011101000111000101010011110101;
	ram[545] = 71'b01011111011001011000100101101011100011111111101000001001111010110111111;
	ram[546] = 71'b01011111010011100011010110011011100101001011101101011110010001010001011;
	ram[547] = 71'b01011111001101101110110101101011001011000000100110110001110011001010011;
	ram[548] = 71'b01011111000111111010111011100010000101100101011001111001011101011011000;
	ram[549] = 71'b01011111000010000111100000001001010110110101011010001001001000111111011;
	ram[550] = 71'b01011110111100010100110011000101101110100000011011100111111010001000000;
	ram[551] = 71'b01011110110110100010100100101100110000010100001111000001001001011110111;
	ram[552] = 71'b01011110110000110000111100101111000101001001000010111101001010010010101;
	ram[553] = 71'b01011110101010111111111011001001100011000101100010000111000011100011000;
	ram[554] = 71'b01011110100101001111011111111001000000100011010011010011110110010001000;
	ram[555] = 71'b01011110011111011111101010111010010100001110111000010111100010010110001;
	ram[556] = 71'b01011110011001110000010100011000101111101110001101101111101100100001000;
	ram[557] = 71'b01011110010100000001101011110100101001001111000111110000110100000100111;
	ram[558] = 71'b01011110001110010011100001101000000001101001011000111001001100000111000;
	ram[559] = 71'b01011110001000100110000101010001111111001101100101111011000110011111001;
	ram[560] = 71'b01011110000010111001000111001101110011110101011010110000110100001011000;
	ram[561] = 71'b01011101111101001100101111001001010101000011001011110100011001101011000;
	ram[562] = 71'b01011101110111100000111101000001011011100010010100001101111011100111001;
	ram[563] = 71'b01011101110001110101101001000011100111010010011000100000110011100111000;
	ram[564] = 71'b01011101101100001011000010101011110111011110110010010110010010101100111;
	ram[565] = 71'b01011101100110100000111010011000100111101000001101001011000010000001000;
	ram[566] = 71'b01011101100000110111010111110110001010011110101011011001101000000000000;
	ram[567] = 71'b01011101011011001110011011000001011010000110010100100011000011011100001;
	ram[568] = 71'b01011101010101100110000011110111010000110101111100100111011001011001101;
	ram[569] = 71'b01011101001111111110010010010100101001010111000010111011111001011000000;
	ram[570] = 71'b01011101001010010110111110101001010000110011000011100000011101101011101;
	ram[571] = 71'b01011101000100110000010000011111110111101111100111111100000111100000001;
	ram[572] = 71'b01011100111111001010000111110101011001101001001001110011000000000000000;
	ram[573] = 71'b01011100111001100100100100100110110010001110101001101011000010100001000;
	ram[574] = 71'b01011100110011111111100110110000111101100001101110000010010110110110111;
	ram[575] = 71'b01011100101110011011000110100101001100101110111110110110011100010111000;
	ram[576] = 71'b01011100101000110111001011101100101110111001000010000000011111000000000;
	ram[577] = 71'b01011100100011010011110110000100100000110100001000111110110110110011101;
	ram[578] = 71'b01011100011101110001000101101001011111100111000110110110000010101101101;
	ram[579] = 71'b01011100011000001110111010011000101000101011001111000111011001000000000;
	ram[580] = 71'b01011100010010101101001100100100110000101000011000111010111100000100101;
	ram[581] = 71'b01011100001101001100000011110101100101100101010010101100110000010001101;
	ram[582] = 71'b01011100000111101011100000001000000101101101101011110100011000000000000;
	ram[583] = 71'b01011100000010001011011001110000000000111110101011111001000000111110101;
	ram[584] = 71'b01011011111100101011111000010100001011100101011000011110101101101110101;
	ram[585] = 71'b01011011110111001100111011110001100100011111110100000101011000000000000;
	ram[586] = 71'b01011011110001101110100100000101001010111110011010010001111000100011000;
	ram[587] = 71'b01011011101100010000110001001011111110100011111110100101011010010111111;
	ram[588] = 71'b01011011100110110011011011011011010001101010000110010001100010011101000;
	ram[589] = 71'b01011011100001010110101010011000011000011111100100111000010011000000000;
	ram[590] = 71'b01011011011011111010011110000000010011011001010010000000010111001111001;
	ram[591] = 71'b01011011010110011110101110101001001111100000100000010101011011111000000;
	ram[592] = 71'b01011011010001000011100011110111100111101111010001011100011101011001000;
	ram[593] = 71'b01011011001011101000111101101000011101001100011000010111111100100010011;
	ram[594] = 71'b01011011000110001110110100010010110111100011000111111111000101111011000;
	ram[595] = 71'b01011011000000110101010110111111111111000110111011111101000111000011101;
	ram[596] = 71'b01011010111011011100010110100001010101100011100011101010101001011011000;
	ram[597] = 71'b01011010110110000011110010110100110110100101111100100000111101100111001;
	ram[598] = 71'b01011010110000101011111011000001111000001010011010000110101000000000000;
	ram[599] = 71'b01011010101011010100011111111011101111101110001001011000000000100101001;
	ram[600] = 71'b01011010100101111101100001100000011001100010001101110110011011001000000;
	ram[601] = 71'b01011010100000100111001110110101011001100110101100111011111101100001011;
	ram[602] = 71'b01011010011011010001011000101111111000101111000111010010100100001000000;
	ram[603] = 71'b01011010010101111011111111001101110011110000011111110001110101111100111;
	ram[604] = 71'b01011010010000100111010001010010111101001001100011111011010110100111000;
	ram[605] = 71'b01011010001011010010111111110110010000101001000001110111011111000110111;
	ram[606] = 71'b01011010000101111111001010110101101011100111110101000011100110010001000;
	ram[607] = 71'b01011010000000101100000001010011001111011110000101111001000011101100001;
	ram[608] = 71'b01011001111011011001010100000111101010011010101101010101111111010001000;
	ram[609] = 71'b01011001110110000111000011010000111010011010011000101110001000101011101;
	ram[610] = 71'b01011001110000110101011101101111010000001001011010100000000100011000000;
	ram[611] = 71'b01011001101011100100010100011101001011111011110111011100101100110001101;
	ram[612] = 71'b01011001100110010011100111011000101100010010001000000000000000000000000;
	ram[613] = 71'b01011001100001000011011110000000000000101110011101100110101111110111000;
	ram[614] = 71'b01011001011011110011111000010000001111110001011010101010010001111011111;
	ram[615] = 71'b01011001010110100100101110100110110100110100011000011010000111101001000;
	ram[616] = 71'b01011001010001010110001000100001000111101111101101110001011001000000000;
	ram[617] = 71'b01011001001100001000000101111100001111110100110100001110011011101100001;
	ram[618] = 71'b01011001000110111010011111010110100001010010011100111001001111111000000;
	ram[619] = 71'b01011001000001101101011100001100011100100100010011001100110110110101000;
	ram[620] = 71'b01011000111100100000111100011011001001101100011111010000100010011000011;
	ram[621] = 71'b01011000110111010100111000100001110101100001101101000111011111101111000;
	ram[622] = 71'b01011000110010001001010000011110100000011000000110000101010100010011011;
	ram[623] = 71'b01011000101100111110001011101100100001000001001101100110100001101010011;
	ram[624] = 71'b01011000100111110011101010001001000000011100101110010001001100010011000;
	ram[625] = 71'b01011000100010101001101011110001000111111100000100000101100110001000000;
	ram[626] = 71'b01011000011101100000001001000101100010001111011110011111001010101000000;
	ram[627] = 71'b01011000011000010111000010000100010000100100100100100000000111001011000;
	ram[628] = 71'b01011000010011001110011110000111001110001010011101010000100000111100011;
	ram[629] = 71'b01011000001110000110011101001011100101001111110101101001101011011001011;
	ram[630] = 71'b01011000001000111110110111110011001011010000110101000001111101110010101;
	ram[631] = 71'b01011000000011110111110101010111000100110011010010011100010101111101000;
	ram[632] = 71'b01010111111110110001001110011001101100100000100101010111100101111011001;
	ram[633] = 71'b01010111111001101011001010010011100010101000110000000000001110100110011;
	ram[634] = 71'b01010111110100100101101001000001110010101001001011001110001000000000000;
	ram[635] = 71'b01010111101111100000100011000111101110110110011010101000010010110000111;
	ram[636] = 71'b01010111101010011011111000100011011010000011011001101001000000000000000;
	ram[637] = 71'b01010111100101010111110000101100001100000101100010111001000110011000000;
	ram[638] = 71'b01010111100000010100001011011111010001010111000001000111001110101000011;
	ram[639] = 71'b01010111011011010001000001100001000110000100101010011001101001011000000;
	ram[640] = 71'b01010111010110001110010010101111101101101101010111110110100011000011111;
	ram[641] = 71'b01010111010001001100001101111001100100001011010010011100101001000011000;
	ram[642] = 71'b01010111001100001010011100110011010010011001011100000011010110010111000;
	ram[643] = 71'b01010111000111001001001110001011000010100010001101100010001010010111001;
	ram[644] = 71'b01010111000010001000100001111110000010011010100011000111001110010010111;
	ram[645] = 71'b01010110111101001000010000110010011100011001011100001101010000111110111;
	ram[646] = 71'b01010110111000001000100001111101000110101011100010011011111101111101000;
	ram[647] = 71'b01010110110011001001001110000100110000001010100011001111100001010001111;
	ram[648] = 71'b01010110101110001010011100011101101011010111000110000111011100001000111;
	ram[649] = 71'b01010110101001001100000101101111001011101000000001001111000110010000001;
	ram[650] = 71'b01010110100100001110010001001100111111110111011001000011000101000111000;
	ram[651] = 71'b01010110011111010000110111011110111111110011100111101010100010010000101;
	ram[652] = 71'b01010110011010010011111000100011010000111110011111110111111011010111000;
	ram[653] = 71'b01010110010101010111011011101100101101000000010001001111000101100001000;
	ram[654] = 71'b01010110010000011011100000111000100100000100000111011101110000100101001;
	ram[655] = 71'b01010110001011100000000000101111110110010111010010101000010111001001000;
	ram[656] = 71'b01010110000110100101000010100100101000100000101001011000001000100111000;
	ram[657] = 71'b01010110000001101010010111101100110010001110011111001001111011110010011;
	ram[658] = 71'b01010101111100110000010110000001011111110100111111010011011100011000000;
	ram[659] = 71'b01010101110111110110101110111000111011010000010010000111010111000001111;
	ram[660] = 71'b01010101110010111101100010010001001011011000100111001110000100101000000;
	ram[661] = 71'b01010101101110000100110111011010111100110010101011001111100101111000000;
	ram[662] = 71'b01010101101001001100100111000001001101101010010101100100011001011011000;
	ram[663] = 71'b01010101100100010100111000010100000111100000110100001011100110100001011;
	ram[664] = 71'b01010101011111011101100011111111001100010101111001100000011100110001000;
	ram[665] = 71'b01010101011010100110101010000000100011110101110010101101001001111101011;
	ram[666] = 71'b01010101010101110000010001100111100011000100011011000010000010110010111;
	ram[667] = 71'b01010101010000111010010011100000100001100011011110101010010011101000101;
	ram[668] = 71'b01010101001100000100110110111010010001100000100100001010100111000011000;
	ram[669] = 71'b01010101000111001111110100100001101110000011111011001010101001101110001;
	ram[670] = 71'b01010101000010011011010011100101000110101010010000000001011110110001111;
	ram[671] = 71'b01010100111101100111001100110001111001111100110101101101100010110101111;
	ram[672] = 71'b01010100111000110011100000000110010000110000111011111001011101111010001;
	ram[673] = 71'b01010100110100000000010100101111100110100001110000011111101010010011000;
	ram[674] = 71'b01010100101111001101100011011100001110111110010000010010110001100100101;
	ram[675] = 71'b01010100101010011011010011011001000010111101110101000001110000010110111;
	ram[676] = 71'b01010100100101101001011101010100111001100011001011010000010000001001011;
	ram[677] = 71'b01010100100000111000000001001101111100010110111011100010100101000000001;
	ram[678] = 71'b01010100011100000111000110010000010000100010101000100011111111101001000;
	ram[679] = 71'b01010100010111010110100101001011100001111010101101110110000011000011101;
	ram[680] = 71'b01010100010010100110100101001011010011010001111101001001101100110100011;
	ram[681] = 71'b01010100001101110110110111110010101100001011001100001001011001111001000;
	ram[682] = 71'b01010100001001000111110010100111001101001010011011110100101101001010101;
	ram[683] = 71'b01010100000100011000111111111111101010101100000100111101001001100011001;
	ram[684] = 71'b01010011111111101010101110010011101010011000111000100001011001000000000;
	ram[685] = 71'b01010011111010111100111101100000100011011001111101111100001000011101000;
	ram[686] = 71'b01010011110110001111011111001100001010111010101011001000010110001010101;
	ram[687] = 71'b01010011110001100010100001101100011111100100010100010100100001100001011;
	ram[688] = 71'b01010011101100110110000100111110111001001001010110010001100000111000000;
	ram[689] = 71'b01010011101000001010000001110101110010000110101111011101001001011110111;
	ram[690] = 71'b01010011100011011110011000001111010110001000111101100100100000101000000;
	ram[691] = 71'b01010011011110110011001000001001110001000101001111000010001100100011011;
	ram[692] = 71'b01010011011010001000011000101101011001001001101111011100110100110101101;
	ram[693] = 71'b01010011010101011110000010101101101110000011001101110100111111100111001;
	ram[694] = 71'b01010011010000110100000110001000111100000100100010010010000001100111111;
	ram[695] = 71'b01010011001100001010101010000110100110101111010000100010010011000000000;
	ram[696] = 71'b01010011000111100001100111011011000001011111100110111001011010001101011;
	ram[697] = 71'b01010011000010111001000101001101001110001011110010000111101100010110001;
	ram[698] = 71'b01010010111110010000110101001001011110100010110101001111011000000000000;
	ram[699] = 71'b01010010111001101001000101011111011000110110001011011101110001111001000;
	ram[700] = 71'b01010010110101000001110110001100010111011100100100111110101110110100111;
	ram[701] = 71'b01010010110000011010111000111110010010010100101110001011100000001000101;
	ram[702] = 71'b01010010101011110100011100000011001010100010111001111100101000111011000;
	ram[703] = 71'b01010010100111001110011000010001001011100011111010101001101111001010001;
	ram[704] = 71'b01010010100010101000110100101101100001110111100011000110111000001011111;
	ram[705] = 71'b01010010011110000011101010001110111011000011010101101010101001001101111;
	ram[706] = 71'b01010010011001011110111000110011100101001111111110000100111111010000001;
	ram[707] = 71'b01010010010100111010100000011001101110101110110000100101110110010001101;
	ram[708] = 71'b01010010010000010110101000000101100001010110101111111010111000011000000;
	ram[709] = 71'b01010010001011110011001000101110101110101011111000111101110101101011101;
	ram[710] = 71'b01010010000111010000000010010011100101011100101110101011000000000000000;
	ram[711] = 71'b01010010000010101101011011110111011101101111101001000101111100101111000;
	ram[712] = 71'b01010001111110001011001110010010111011111011001100001100111111001111000;
	ram[713] = 71'b01010001111001101001011001100100001111001011000100100101000000000000000;
	ram[714] = 71'b01010001110101000111111101101001100110110011100011110001011001001000000;
	ram[715] = 71'b01010001110000100110111010100001010010010001011111110111010010101101000;
	ram[716] = 71'b01010001101100000110010111001101010111000101010010001001011101001101011;
	ram[717] = 71'b01010001100111100110001100100111101101110011111101101000101000011111000;
	ram[718] = 71'b01010001100011000110100001110001111011000110011001001001001111011000000;
	ram[719] = 71'b01010001011110100111001000100011010100111100011110111110111110110100011;
	ram[720] = 71'b01010001011010001000001111000000100100011101010000111111111001111110101;
	ram[721] = 71'b01010001010101101001101110000100100101010000100100010111111001000000001;
	ram[722] = 71'b01010001010001001011100101101101100111110101101110011100000011011000111;
	ram[723] = 71'b01010001001100101101111100111011111110111010000111111100011000000000000;
	ram[724] = 71'b01010001001000010000101100101011011000001011111000011100110011110110011;
	ram[725] = 71'b01010001000011110011110100111010000100100111001011011001110101000000000;
	ram[726] = 71'b01010000111111010111010101100110010101010000101011010011111111100010111;
	ram[727] = 71'b01010000111010111011001110101110011011010101100001010011011101000000000;
	ram[728] = 71'b01010000110110011111100111010001011000000101101101001000101011011000000;
	ram[729] = 71'b01010000110010000100011000001100001100010100001011000010011000101001000;
	ram[730] = 71'b01010000101101101001100001011101001001101010110010010100100110110101000;
	ram[731] = 71'b01010000101001001111000011000010100001111011110110111101110010001000000;
	ram[732] = 71'b01010000100100110101000011111010010101100010111000011111111111100010001;
	ram[733] = 71'b01010000100000011011010110000011001001001101110100101101101100111011111;
	ram[734] = 71'b01010000011100000010000111011010011011111000101001100111001000000000000;
	ram[735] = 71'b01010000010111101001010000111110110001011001111110010101101010110011011;
	ram[736] = 71'b01010000010011010000111001101101001001101011100101001110001001000101001;
	ram[737] = 71'b01010000001110111000110011100110001100010010101011000010111000000000000;
	ram[738] = 71'b01010000001010100001001100100101010110100111100011011000010010001101000;
	ram[739] = 71'b01010000000110001001111101101010001110001100011101010010111000101011000;
	ram[740] = 71'b01010000000001110011000110110011000110000110000001110000110001001000000;
	ram[741] = 71'b01001111111101011100100111111110010001100001010001101001000001001000000;
	ram[742] = 71'b01001111111001000110100001001010000011110011100101001111100100101011000;
	ram[743] = 71'b01001111110100110000111001010001101100100110010001001110100100101010011;
	ram[744] = 71'b01001111110000011011100010011001010111000001011101010111111111001010001;
	ram[745] = 71'b01001111101100000110101010011000111111000110100011010111010010100101000;
	ram[746] = 71'b01001111100111110010001010010001111100100100000010010101011001111111101;
	ram[747] = 71'b01001111100011011110000010000010100011011100010011110101111110011001000;
	ram[748] = 71'b01001111011111001010011000100100110011110000101001110001110011110001000;
	ram[749] = 71'b01001111011010110110111111111111011010000110000100100011100011110101011;
	ram[750] = 71'b01001111010110100100000110000111110010100110101101000001110010110010111;
	ram[751] = 71'b01001111010010010001100100000000100110000010111011000100101101110000101;
	ram[752] = 71'b01001111001101111111011001101000001001001001111100111110101111111001101;
	ram[753] = 71'b01001111001001101101100110111100110000110011010011010100101110000101111;
	ram[754] = 71'b01001111000101011100001011111100110001111110110000100001111111110010011;
	ram[755] = 71'b01001111000001001011001000100110100001110100011000011100101001010011001;
	ram[756] = 71'b01001110111100111010100011110010000001110101100100000001110000001101000;
	ram[757] = 71'b01001110111000101010001111101001111111000000111110110001100111011000000;
	ram[758] = 71'b01001110110100011010011001111111110111100100011001111101001011000010001;
	ram[759] = 71'b01001110110000001010111011111000010100111011000111100101000011000000000;
	ram[760] = 71'b01001110101011111011110101010001101100111001101100110110110000000000001;
	ram[761] = 71'b01001110100111101101000110001010010101011100111101101000110110011000000;
	ram[762] = 71'b01001110100011011110101110100000100100101001111011111111010010111001001;
	ram[763] = 71'b01001110011111010000101110010010110000101101110111101111110001000000000;
	ram[764] = 71'b01001110011011000011001100010110111101110010110000000101101000000101000;
	ram[765] = 71'b01001110010110110101111010111011110110111110011111100011111101000110101;
	ram[766] = 71'b01001110010010101001000111101110111110110011111001100010000111001111011;
	ram[767] = 71'b01001110001110011100101011110110111110001111101110100001110100010100011;
	ram[768] = 71'b01001110001010010000100111010010001100001011011100100001001010010101101;
	ram[769] = 71'b01001110000110000100111001111110111111101000101100011111100001001110001;
	ram[770] = 71'b01001110000001111001100011111011101111110001010010000010000011100101111;
	ram[771] = 71'b01001101111101101110100101000110110011110111001010111000010000111101111;
	ram[772] = 71'b01001101111001100011111101011110100011010100011110100000100001010110001;
	ram[773] = 71'b01001101110101011001101101000001010101101011011101101100101010001101101;
	ram[774] = 71'b01001101110001001111110011101101100010100110100010000110100100111100011;
	ram[775] = 71'b01001101101101000110011000010110100011101011001001001101011001001000000;
	ram[776] = 71'b01001101101000111101001101010000011101101011101100110001100011000111000;
	ram[777] = 71'b01001101100100110100100000000011011100110000111110111111011110110000011;
	ram[778] = 71'b01001101100000101100000011000100100100000110011011100000011111110011001;
	ram[779] = 71'b01001101011100100100000011111011000010000000100010010111100001010101000;
	ram[780] = 71'b01001101011000011100011011110000101100001110000001000000101010000110101;
	ram[781] = 71'b01001101010100010101001010100011111011010101010001001110100011100001000;
	ram[782] = 71'b01001101010000001110010000010011001000000100110010000110101000110001001;
	ram[783] = 71'b01001101001100000111100110001001100101010010111010000001011001011010001;
	ram[784] = 71'b01001101001000000001011001101100000111011000000110111011101001011000000;
	ram[785] = 71'b01001101000011111011100100000101110010000000011000110000110101010111001;
	ram[786] = 71'b01001100111111110110001100000111010110010001101011011000011101111011001;
	ram[787] = 71'b01001100111011110001000100001010001110011110001101010111111100001101000;
	ram[788] = 71'b01001100110111101100010010111111011011010011010001111011010100111010101;
	ram[789] = 71'b01001100110011100111111000100101010110010111110001010011011000001001000;
	ram[790] = 71'b01001100101111100011110100111010011001011010100101101010101101010001001;
	ram[791] = 71'b01001100101011100000000111111100111110010010101010101010110010000001000;
	ram[792] = 71'b01001100100111011100111000011100011011000001010101000001111101100111000;
	ram[793] = 71'b01001100100011011001111000110101000010011000111110101011101101000100011;
	ram[794] = 71'b01001100011111010111001111110110011001111011110100101101111011011101000;
	ram[795] = 71'b01001100011011010101000100001111001010010111011000000111010001111000000;
	ram[796] = 71'b01001100010111010011001000011101000010010000110111000110111111010001111;
	ram[797] = 71'b01001100010011010001100011001110111001110011011100001001111111001000000;
	ram[798] = 71'b01001100001111010000011011010010101100100010010101000010101010111000000;
	ram[799] = 71'b01001100001011001111100011000111100100100010010111011110101101110101101;
	ram[800] = 71'b01001100000111001111000001011011101100110001001100001110001000000000000;
	ram[801] = 71'b01001100000011001110111100111100010011110001001101010010101010010111000;
	ram[802] = 71'b01001011111111001111001000001001111110110011101101010100101011010010101;
	ram[803] = 71'b01001011111011001111110000100000100001000010110111100110001111010101111;
	ram[804] = 71'b01001011110111010000101000100001011100011000000011011011110101011001000;
	ram[805] = 71'b01001011110011010001110110111001110000101111100101010110100000000000111;
	ram[806] = 71'b01001011101111010011100010010101100001111111101100010111010000001011111;
	ram[807] = 71'b01001011101011010101011101010111101100101110010101011111101101000000000;
	ram[808] = 71'b01001011100111010111101110101100100100000011100101111001111000100101011;
	ram[809] = 71'b01001011100011011010011100111111011111001110000111001100000011101000001;
	ram[810] = 71'b01001011011111011101011010110100110101001101010111100011101000000000000;
	ram[811] = 71'b01001011011011100000101110111000001100011110101001101000110101010100001;
	ram[812] = 71'b01001011010111100100011001001000000001011111110111000000110000101000000;
	ram[813] = 71'b01001011010011101000100000001110110000001110101110100111101101111101000;
	ram[814] = 71'b01001011001111101100110110110010100111101111011010011101111010111100001;
	ram[815] = 71'b01001011001011110001100011011110010011001010000001101000100111000101000;
	ram[816] = 71'b01001011000111110110100110010000001111011011111100010011100101101101101;
	ram[817] = 71'b01001011000011111011111111000110111001101010011001010010110101101001000;
	ram[818] = 71'b01001011000000000001101110000000101111000010011101101000000110000110001;
	ram[819] = 71'b01001010111100000111110010111100001100111001000100001000011101001001000;
	ram[820] = 71'b01001010111000001110001101110111110000101010111101000001111111011101101;
	ram[821] = 71'b01001010110100010100111110110001110111111100101101100001011001100101000;
	ram[822] = 71'b01001010110000011100000101101001000000011010101111010111101010011100001;
	ram[823] = 71'b01001010101100100011011011110001111100110001111101101111111101110011001;
	ram[824] = 71'b01001010101000101011001110011110101111111100000110101111000100101000000;
	ram[825] = 71'b01001010100100110011010111000011111110000101100010110101000000011100001;
	ram[826] = 71'b01001010100000111011101110110111000110011101001100110000111110111101111;
	ram[827] = 71'b01001010011101000100100011001000110011111011111000000000000000000000000;
	ram[828] = 71'b01001010011001001101100110100101110101101101101000111110100101001001000;
	ram[829] = 71'b01001010010101010110111111110101101001001111000011001010100000101011000;
	ram[830] = 71'b01001010010001100000110101011110110001011001100101111000111000001000101;
	ram[831] = 71'b01001010001101101010111010001111010101110000101101100000100011101101101;
	ram[832] = 71'b01001010001001110101010100101110001000000110101010101011110111010101111;
	ram[833] = 71'b01001010000110000000000100111001100111011010010110111101111110011110011;
	ram[834] = 71'b01001010000010001011001010110000010010110010011011101110011110011011001;
	ram[835] = 71'b01001001111110010110100110010000101001011101010001101111010010100011001;
	ram[836] = 71'b01001001111010100010010111011001001010110001000000110010101001110110011;
	ram[837] = 71'b01001001110110101110010111100001110111111101001110110001101010110111000;
	ram[838] = 71'b01001001110010111010110011110110011011100100111101001110100111101000000;
	ram[839] = 71'b01001001101111000111011111001000100111011000001110000110100101000100011;
	ram[840] = 71'b01001001101011010100100110100011001100000100111011111100010110101011101;
	ram[841] = 71'b01001001100111100001111100111000110101101010111100011000111000000000000;
	ram[842] = 71'b01001001100011101111101000101110000101011000100011111011001001010100101;
	ram[843] = 71'b01001001011111111101101010000001011011010110110001101101001011011000000;
	ram[844] = 71'b01001001011100001100000000110001010111110110010000110100000111010000101;
	ram[845] = 71'b01001001011000011010101100111100011011001111010111110110011000000000000;
	ram[846] = 71'b01001001010100101001101110100001000110000010001000100001110101011111101;
	ram[847] = 71'b01001001010000111001000101011101111000110110001111010010000000111000000;
	ram[848] = 71'b01001001001101001000101011001101010101000010001010010010001010101000000;
	ram[849] = 71'b01001001001001011000100110010010010111100010001000000101111101010111000;
	ram[850] = 71'b01001001000101101000111101001111000011111110111001010001111010011010011;
	ram[851] = 71'b01001001000001111001100010111010100111101101000000001011001110000011001;
	ram[852] = 71'b01001000111110001010011101110111010100111001110100110010100111010111001;
	ram[853] = 71'b01001000111010011011101110000011101100110111110110010000001111110110011;
	ram[854] = 71'b01001000110110101101001100111011100111011111000011010101001011100111000;
	ram[855] = 71'b01001000110010111111000111100011000111100101101000010101111101101000000;
	ram[856] = 71'b01001000101111010001010000110011101001111111001100111110111111001000011;
	ram[857] = 71'b01001000101011100011110101110000011000101111100111001001011111011011101;
	ram[858] = 71'b01001000100111110110101001010011101001110111001010001100001000000000000;
	ram[859] = 71'b01001000100100001001110001111110001100010101010010110101100001011100101;
	ram[860] = 71'b01001000100000011101001111101110100010001110101011111001110000011000000;
	ram[861] = 71'b01001000011100110000111100000010000111101011101010111111001100111000000;
	ram[862] = 71'b01001000011001000101000011111001111001010001010101101100000111001101111;
	ram[863] = 71'b01001000010101011001011010010010011011011011000001111110000000001011011;
	ram[864] = 71'b01001000010001101110000101101011010110101100100100100110010110111101001;
	ram[865] = 71'b01001000001110000011001100100011011011010000100111000111010011001001000;
	ram[866] = 71'b01001000001010011000011011011000100011001100101001000000101111100010011;
	ram[867] = 71'b01001000000110101110000101101001111010000000110001011011010000100110111;
	ram[868] = 71'b01001000000011000100000100110101110101000111111100101010011100001011101;
	ram[869] = 71'b01000111111111011010010010011011100010010101110110100101110111001000000;
	ram[870] = 71'b01000111111011110000110100111001010110001101010110111100111001001011101;
	ram[871] = 71'b01000111111000000111101100001101110100000000001000010010101101000000000;
	ram[872] = 71'b01000111110100011110111000010111011111000111010110100010011001001110101;
	ram[873] = 71'b01000111110000110110011001010100111011000011101110100101101110101000000;
	ram[874] = 71'b01000111101101001110001000100110011100001011111110001001001001111000000;
	ram[875] = 71'b01000111101001100110010011000111010010101111110000101010111011110010111;
	ram[876] = 71'b01000111100101111110101011111001110001111110101001011100011110000001011;
	ram[877] = 71'b01000111100010010111011001011010101101000101110010100111101000010100001;
	ram[878] = 71'b01000111011110110000010101001011010000100110001101010011111000000000000;
	ram[879] = 71'b01000111011011001001101100000100111101101000000110011110011110000001000;
	ram[880] = 71'b01000111010111100011010001001011110111010000111111001111011100000101101;
	ram[881] = 71'b01000111010011111101001010111011111001011001100010100110110010101101000;
	ram[882] = 71'b01000111010000010111011001010011101000011111110000111010010111011000001;
	ram[883] = 71'b01000111001100110001111100010001101001001001000111110111000101110101000;
	ram[884] = 71'b01000111001001001100101101011000011011101011011011110000101000101000000;
	ram[885] = 71'b01000111000101100111111001011110111011011100111001011101101000110110001;
	ram[886] = 71'b01000111000010000011010011101011110010011101001000011001001100100001111;
	ram[887] = 71'b01000110111110011111000010011001101010000011011100101110110111001101111;
	ram[888] = 71'b01000110111010111010111111001011111010001010011101011101111000000000000;
	ram[889] = 71'b01000110110111010111010110110111110000001011010011110100101111101000000;
	ram[890] = 71'b01000110110011110011111100100101100100110000110010010110010110001101001;
	ram[891] = 71'b01000110110000010000110110101111001010100010110100001011000000000000000;
	ram[892] = 71'b01000110101100101110000101010011000111000011101100001100001111101011001;
	ram[893] = 71'b01000110101001001011100001110101110111010111111100111100001101110101011;
	ram[894] = 71'b01000110100101101001011001001010100000000110010111111111000000000000000;
	ram[895] = 71'b01000110100010000111011110011011100011100110110111110000101111010111000;
	ram[896] = 71'b01000110011110100101110001101000010000110110100011000010101000010100101;
	ram[897] = 71'b01000110011011000100011111100010011010101100001110001000010110101001111;
	ram[898] = 71'b01000110010111100011011011010101110101110000110011101000010111110001000;
	ram[899] = 71'b01000110010100000010101011011010100111111001001101001001110111011000111;
	ram[900] = 71'b01000110010000100010001111101111010111011100110001000110100111010111000;
	ram[901] = 71'b01000110001101000010001000010010101010111010001100110111001110000010111;
	ram[902] = 71'b01000110001001100010001110101010111010111010011011010101010110010000001;
	ram[903] = 71'b01000110000110000010101001001111010111001110101001010010101010000100101;
	ram[904] = 71'b01000110000010100011010111111110100110101000100111001001111011110000011;
	ram[905] = 71'b01000101111111000100011010110111010000000001011010111011111011101000011;
	ram[906] = 71'b01000101111011100101101011100000100010100100110100111010011011111000000;
	ram[907] = 71'b01000101111000000111010000010000111000001110101100100000011100100111111;
	ram[908] = 71'b01000101110100101001001001000110111000001011000111000001111000001000000;
	ram[909] = 71'b01000101110001001011010110000001001001101101011110000000000001111110011;
	ram[910] = 71'b01000101101101101101110000100111110010010101111000100101011100101001011;
	ram[911] = 71'b01000101101010010000011111010000010110011001001110001100010000110000101;
	ram[912] = 71'b01000101100110110011100001111001011101011101110011111010101001100111001;
	ram[913] = 71'b01000101100011010110110010001011110101101001000011001000101111000011000;
	ram[914] = 71'b01000101011111111010010110011100011011001011001001001111101100010111101;
	ram[915] = 71'b01000101011100011110001110101001110101111101010100001111000100110011000;
	ram[916] = 71'b01000101011001000010011010110010101110000000000011111011111011011111001;
	ram[917] = 71'b01000101010101100110110100100000100111010100010001001110111011000100101;
	ram[918] = 71'b01000101010010001011100010000111101000111011110001001100111010011001011;
	ram[919] = 71'b01000101001110110000100011100110011011001001111000110111010100001010011;
	ram[920] = 71'b01000101001011010101110010100111001010010010001100011000010010001000000;
	ram[921] = 71'b01000101000111111011011011110001100100010111101111100001000000000000000;
	ram[922] = 71'b01000101000100100001010010011011100111000111001010100101011011001100101;
	ram[923] = 71'b01000101000001000111010110100100100011000101100011011000001101100100011;
	ram[924] = 71'b01000100111101101101101110011111001111111000011000001100010000001000011;
	ram[925] = 71'b01000100111010010100011010001010010110011000100000011001111011111000101;
	ram[926] = 71'b01000100110110111011011001100100011111100110000001111000111101100000001;
	ram[927] = 71'b01000100110011100010100110011001010101010111011000100011011000101011000;
	ram[928] = 71'b01000100110000001010001101001101101100101001111001000010011011110111000;
	ram[929] = 71'b01000100101100110001111011000111111000100101111111010001111101100011000;
	ram[930] = 71'b01000100101001011010000010111110111000110000000000100110011111111100001;
	ram[931] = 71'b01000100100110000010011000001100011010000101000000010010001001010010101;
	ram[932] = 71'b01000100100010101011000001000001101011000001011010010000010110000000011;
	ram[933] = 71'b01000100011111010011110111001011100101000100010100001100001001001101000;
	ram[934] = 71'b01000100011011111101000000111010111100011111010000111110100101110100011;
	ram[935] = 71'b01000100011000100110011110001110011011001010010011000110110011110111000;
	ram[936] = 71'b01000100010101010000001111000100101011000100101000001110101011111011011;
	ram[937] = 71'b01000100010001111010001101001011011010100010110010010111001101011101001;
	ram[938] = 71'b01000100001110100100011110110010101001101101010011001100101000110010001;
	ram[939] = 71'b01000100001011001110111101101000100001001100111111111110100001101101000;
	ram[940] = 71'b01000100000111111001110110001100111011101111011101111100000001001011000;
	ram[941] = 71'b01000100000100100100111011111101101101100100001000010111100110011111011;
	ram[942] = 71'b01000100000001010000001110111010001000010101111000000000110110001100001;
	ram[943] = 71'b01000011111101111011110101010001001011010011010100001001011001011100001;
	ram[944] = 71'b01000011111010100111101111000001100001001100000100001000111110001111011;
	ram[945] = 71'b01000011110111010011111100001001110100110110110111100111000001100110111;
	ram[946] = 71'b01000011110100000000010110011001101010101100010100110111110110011000000;
	ram[947] = 71'b01000011110000101101000011111111001110010000100001110011011101010101011;
	ram[948] = 71'b01000011101101011001111110101010011110000001000000100001001000101000011;
	ram[949] = 71'b01000011101010000111001100101001001011110000011001000011111010010111101;
	ram[950] = 71'b01000011100110110100101101111010000010110011001000111111010111111110001;
	ram[951] = 71'b01000011100011100010011100001101101000101001010001010010101011001111000;
	ram[952] = 71'b01000011100000010000011101110001001000100010100111000110000101110110101;
	ram[953] = 71'b01000011011100111110110010100011001110000101111111001010010001111111000;
	ram[954] = 71'b01000011011001101101010100010101000101101110001111110111001000000000000;
	ram[955] = 71'b01000011010110011100001001010011010100010000000000010000001011001000000;
	ram[956] = 71'b01000011010011001011010001011100100101100100011001101100111110000101000;
	ram[957] = 71'b01000011001111111010100110100010101100111001011111010100101111011110001;
	ram[958] = 71'b01000011001100101010001110110001101000110000001110000111010001001101000;
	ram[959] = 71'b01000011001001011010001010001000000101010100000001011101001010111111101;
	ram[960] = 71'b01000011000110001010010010011000011100011110100001011001010010001100001;
	ram[961] = 71'b01000011000010111010100111100010000000111101100000100111001110011111000;
	ram[962] = 71'b01000010111111101011010101111011110111001101001101110101100000001111000;
	ram[963] = 71'b01000010111100011100010001001100101101010011001001000101100110011111111;
	ram[964] = 71'b01000010111001001101011001010011110110000111101110101111101111111100001;
	ram[965] = 71'b01000010110101111110111010100111001001110111101100001001110001111011000;
	ram[966] = 71'b01000010110010110000100010100011011101011011100111000001100110111010011;
	ram[967] = 71'b01000010101111100010100011101001010101101001111010101001011011101001011;
	ram[968] = 71'b01000010101100010100110001100001100000010111111001111100011101111000000;
	ram[969] = 71'b01000010101001000111001100001011010000101111001000001101111011101011000;
	ram[970] = 71'b01000010100101111001111111111010100000010111011000010001111010001001011;
	ram[971] = 71'b01000010100010101101000000011001001001011100010111110110011010011000001;
	ram[972] = 71'b01000010011111100000001101100110011111010010001111010111111000000000000;
	ram[973] = 71'b01000010011100010011101101101011100010100011110110110001011111011100001;
	ram[974] = 71'b01000010011001000111100000100111000000110100100100100000001101101000000;
	ram[975] = 71'b01000010010101111011100000001110010011100110111100000000100001000000000;
	ram[976] = 71'b01000010010010101111110010101001110101111110001001100001100000011111000;
	ram[977] = 71'b01000010001111100100010001101111011010110001101110100100110111001001101;
	ram[978] = 71'b01000010001100011001000011100111000100000010111100000000101010000111000;
	ram[979] = 71'b01000010001001001110001000001111011111110010001110011111110111001111001;
	ram[980] = 71'b01000010000110000011011001011111000110110001101111000011011011001011101;
	ram[981] = 71'b01000010000010111000111101011101010101100111000111100001111000100111011;
	ram[982] = 71'b01000001111111101110101110000000111110010001010111110111110010110001000;
	ram[983] = 71'b01000001111100100100110001010001000100011100010001000110001001110111011;
	ram[984] = 71'b01000001111001011011000111001100010110100101001111011001100110001011000;
	ram[985] = 71'b01000001110110010001101001101010001100011001110000010111100110001101000;
	ram[986] = 71'b01000001110011001000011000101001111001111100101001111110010010110001111;
	ram[987] = 71'b01000001101111111111011010010001110001001111011110110101101110000011000;
	ram[988] = 71'b01000001101100110110101110100000100001000101101001011110010111100111111;
	ram[989] = 71'b01000001101001101110010101010100111000011001011110111110000110111101000;
	ram[990] = 71'b01000001100110100110001000100111001101011111111100010111100100010011000;
	ram[991] = 71'b01000001100011011110001000010110110100101100101010110010010010001111011;
	ram[992] = 71'b01000001100000010110011010101001000010001111011000111111010100101001000;
	ram[993] = 71'b01000001011101001110111111011100100101011000010101010000001011001011011;
	ram[994] = 71'b01000001011010000111110000101010100110010011001010011100111001110101101;
	ram[995] = 71'b01000001010111000000110100010111110100010101001011100010111101111111001;
	ram[996] = 71'b01000001010011111010000100011101110000100000100111111000000101011111000;
	ram[997] = 71'b01000001010000110011100111000000110001100110111111011100001011000101101;
	ram[998] = 71'b01000001001101101101010101111010110001011110000010000110101111100110101;
	ram[999] = 71'b01000001001010100111010111001111101110010110011111000111101111010010111;
	ram[1000] = 71'b01000001000111100001100100111001111010110110100011001010011101110001000;
	ram[1001] = 71'b01000001000100011100000100111100111100110001001110101110110000001111111;
	ram[1002] = 71'b01000001000001010110110111010111100100001001001101100000100100001111000;
	ram[1003] = 71'b01000000111110010001110110000100101000101000100101101100101111011111000;
	ram[1004] = 71'b01000000111011001101000111000111001011011100111101111001000000000000000;
	ram[1005] = 71'b01000000111000001000100100011010011100111000111000100001011011100011011;
	ram[1006] = 71'b01000000110101000100010100000001000101110100001001011111000101000000000;
	ram[1007] = 71'b01000000110010000000001111110110101111000110101100100001001001110111000;
	ram[1008] = 71'b01000000101110111100011101111101101001010101100100000010100110100011000;
	ram[1009] = 71'b01000000101011111000111000010001110101111011000010010111011000111011111;
	ram[1010] = 71'b01000000101000110101100100110101001101001100011001011101010100111101000;
	ram[1011] = 71'b01000000100101110010011101100100001001000011001111101100100001000011000;
	ram[1012] = 71'b01000000100010101111101000100000001001101000000111011001000001001000000;
	ram[1013] = 71'b01000000011111101100111111100110000001010000111000101100001010110001011;
	ram[1014] = 71'b01000000011100101010101000110110110111111100010110110110000110001000000;
	ram[1015] = 71'b01000000011001101000100100010001011110110100111001111010001010111100111;
	ram[1016] = 71'b01000000010110100110101011110011001100110110000101001010100101010010011;
	ram[1017] = 71'b01000000010011100100111111011011010111100111000011100001000000000000000;
	ram[1018] = 71'b01000000010000100011100101001010010110111100100011000001111001110000111;
	ram[1019] = 71'b01000000001101100010010110111110000110001110101101011101111100100101111;
	ram[1020] = 71'b01000000001010100001011010110110100101010001100010010101001011011011001;
	ram[1021] = 71'b01000000000111100000110000110010100101101111100111101011101110001111101;
	ram[1022] = 71'b01000000000100100000010010110000100111011001001011000001001000000001000;
	ram[1023] = 71'b01000000000001100000000000110000000000001000000000000000000000000000000;
end
endmodule
`default_nettype wire