// load_tableをノンブロッキング代入すべきかは要調査。

`default_nettype none
module finv_load_const_table (
    input wire [9:0] addr,
    output wire [57:0] cst,
    input wire clk,
	input wire rstn);

(* RAM_STYLE="BLOCK" *) reg [57:0] ram [1023:0];
//always @(posedge clk)
//    cst <= ram[addr];
assign cst = ram[addr];
initial begin
	ram[0] = 58'b1111111111111111111111000000000111111111110000000000000000;
	ram[1] = 58'b1111111111000000000011000000000100000001001111100111000000;
	ram[2] = 58'b1111111110000000001110111110100000010110101010101110000000;
	ram[3] = 58'b1111111101000000100010111001111100101010000010101111101101;
	ram[4] = 58'b1111111100000000111110110000111011111100011011010100111100;
	ram[5] = 58'b1111111011000001100010100001111100100111110110100111000011;
	ram[6] = 58'b1111111010000010001110001011100011011011111110100110100000;
	ram[7] = 58'b1111111001000011000001101100001111100010000100101011111001;
	ram[8] = 58'b1111111000000011111101000010100101011000100111111111100000;
	ram[9] = 58'b1111110111000101000000001101000111110110000001000101011111;
	ram[10] = 58'b1111110110000110001011001010011000001001000010001100011000;
	ram[11] = 58'b1111110101000111011101111000111010110101101001110100000000;
	ram[12] = 58'b1111110100001000111000010111010100110110011011010101010000;
	ram[13] = 58'b1111110011001010011010100100001000011110111101011011001100;
	ram[14] = 58'b1111110010001100000100011101111011010111001010110101010010;
	ram[15] = 58'b1111110001001101110110000011010010011110001101000101010001;
	ram[16] = 58'b1111110000001111101111010010110010001010101001001101110000;
	ram[17] = 58'b1111101111010001110000001011000000001000011110001100110111;
	ram[18] = 58'b1111101110010011111000101010100100010111100000110010001110;
	ram[19] = 58'b1111101101010110001000110000000010010011010010111100010100;
	ram[20] = 58'b1111101100011000100000011010000010100111100110011011000000;
	ram[21] = 58'b1111101011011010111111100111001011011001100111001100000000;
	ram[22] = 58'b1111101010011101100110010110000100000011000110010011101000;
	ram[23] = 58'b1111101001100000010100100101010100010011011101111010100100;
	ram[24] = 58'b1111101000100011001010010011100011010001001100010101101000;
	ram[25] = 58'b1111100111100110000111011111011011010011101010101001101111;
	ram[26] = 58'b1111100110101001001100000111100011001101101101110101100000;
	ram[27] = 58'b1111100101101100011000001010100101000010110001001100111101;
	ram[28] = 58'b1111100100101111101011100111001010001100111010000100000000;
	ram[29] = 58'b1111100011110011000110011011111011011101000100011000001100;
	ram[30] = 58'b1111100010110110101000100111100010110111011110100001000010;
	ram[31] = 58'b1111100001111010010010001000101011110011001111111111000100;
	ram[32] = 58'b1111100000111110000010111110000000000000000000000000000000;
	ram[33] = 58'b1111100000000001111011000110001010100000001001111010111111;
	ram[34] = 58'b1111011111000101111010011111110110101010101011100010101110;
	ram[35] = 58'b1111011110001010000001001001110000001010111110111011010000;
	ram[36] = 58'b1111011101001110001111000010100011000000110100001111110000;
	ram[37] = 58'b1111011100010010100100001000111011100000001011101000010011;
	ram[38] = 58'b1111011011010111000000011011100101010011100101011010100000;
	ram[39] = 58'b1111011010011011100011111001001110010101000000100001000000;
	ram[40] = 58'b1111011001100000001110100000100011110100101000100111011000;
	ram[41] = 58'b1111011000100101000000010000010010011001000010010111111100;
	ram[42] = 58'b1111010111101001111001000111001000110111101001000110000000;
	ram[43] = 58'b1111010110101110111001000011110100011110100110100100110100;
	ram[44] = 58'b1111010101110100000000000101000011101101001101000000000000;
	ram[45] = 58'b1111010100111001001110001001100101010110001110100100101100;
	ram[46] = 58'b1111010011111110100011010000001001011101000100001001110010;
	ram[47] = 58'b1111010011000011111111010111011101100000110010100110000001;
	ram[48] = 58'b1111010010001001100010011110010011001000011110011101000000;
	ram[49] = 58'b1111010001001111001100100011011000011001110011000111000000;
	ram[50] = 58'b1111010000010100111101100101011110100100110101000101111000;
	ram[51] = 58'b1111001111011010110101100011010101010010100100000100011101;
	ram[52] = 58'b1111001110100000110100011011101111010101101001100011001100;
	ram[53] = 58'b1111001101100110111010001101011011111111111001000010001100;
	ram[54] = 58'b1111001100101101000110110111001100101111101110011001101000;
	ram[55] = 58'b1111001011110011011010010111110100010010111000000110100100;
	ram[56] = 58'b1111001010111001110100101110000011110000001000001101001000;
	ram[57] = 58'b1111001010000000010101111000101101011101011111101101001111;
	ram[58] = 58'b1111001001000110111101110110100100000011010110010110000000;
	ram[59] = 58'b1111001000001101101100100110011011011000110010101100000101;
	ram[60] = 58'b1111000111010100100010000111000100110001101011110001000000;
	ram[61] = 58'b1111000110011011011110010111010101100101110100011111011011;
	ram[62] = 58'b1111000101100010100001010101111111101101011010001000100000;
	ram[63] = 58'b1111000100101001101011000001111000000111101111100100000000;
	ram[64] = 58'b1111000011110000111011011001110011001001100100101111000000;
	ram[65] = 58'b1111000010111000010010011100100100011101010010111111000000;
	ram[66] = 58'b1111000001111111110000001001000010110011011011101001101110;
	ram[67] = 58'b1111000001000111010100011110000000100001100110001000010101;
	ram[68] = 58'b1111000000001110111111011010010100111011011000111111000000;
	ram[69] = 58'b1110111111010110110000111100110100110001101101110110101011;
	ram[70] = 58'b1110111110011110101001000100010110111110110000111110101010;
	ram[71] = 58'b1110111101100110100111101111110000110110001101001101100001;
	ram[72] = 58'b1110111100101110101100111101111000111000111000100010111000;
	ram[73] = 58'b1110111011110110111000101101100101111000110001011101111111;
	ram[74] = 58'b1110111010111111001010111101101110111000111010000000110110;
	ram[75] = 58'b1110111010000111100011101101001010010001101101110100000000;
	ram[76] = 58'b1110111001010000000010111010110001011111010100101101010000;
	ram[77] = 58'b1110111000011000101000100101011011011011110101001011001100;
	ram[78] = 58'b1110110111100001010100101011111111010010010011100101100010;
	ram[79] = 58'b1110110110101010000111001101010110010101011011011000000100;
	ram[80] = 58'b1110110101110011000000001000011000010001101000111011000000;
	ram[81] = 58'b1110110100111011111111011011111110111010101000011001110000;
	ram[82] = 58'b1110110100000101000101000111000011011001000111111000000000;
	ram[83] = 58'b1110110011001110010001001000011101001111111010011001010000;
	ram[84] = 58'b1110110010010111100011011111000111111110111001101010110000;
	ram[85] = 58'b1110110001100000111100001001111101011111101101001111101100;
	ram[86] = 58'b1110110000101010011011000111110110000110000111110111101000;
	ram[87] = 58'b1110101111110100000000010111101110000010001011111110010000;
	ram[88] = 58'b1110101110111101101011111000011110000111111111100110100000;
	ram[89] = 58'b1110101110000111011101101001000011000111010011110110111100;
	ram[90] = 58'b1110101101010001010101101000010110010100001111011111011000;
	ram[91] = 58'b1110101100011011010011110101010100000011010001110001011101;
	ram[92] = 58'b1110101011100101011000001110110111111101101111111001100100;
	ram[93] = 58'b1110101010101111100010110011111101111100101000101100000000;
	ram[94] = 58'b1110101001111001110011100011100001001101111011111110100010;
	ram[95] = 58'b1110101001000100001010011100011111000100011001100100010001;
	ram[96] = 58'b1110101000001110100111011101110011001101000101000110100000;
	ram[97] = 58'b1110100111011001001010100110011011011001011100000000000000;
	ram[98] = 58'b1110100110100011110011110101010011110101010100000011011110;
	ram[99] = 58'b1110100101101110100011001001011001110110010011001000010100;
	ram[100] = 58'b1110100100111001011000100001101011111011011010010111000000;
	ram[101] = 58'b1110100100000100010011111101000110111110001010000000001100;
	ram[102] = 58'b1110100011001111010101011010101001000001011011101010000000;
	ram[103] = 58'b1110100010011010011100111001010000010111000110110110100100;
	ram[104] = 58'b1110100001100101101010010111111010100101111001110101011000;
	ram[105] = 58'b1110100000110000111101110101101000010001100100110001101111;
	ram[106] = 58'b1110011111111100010111010001010111011110011001011000010110;
	ram[107] = 58'b1110011111000111110110101010000110011111100011101101000000;
	ram[108] = 58'b1110011110010011011011111110110101101010110001101111010100;
	ram[109] = 58'b1110011101011111000111001110100100101010010110101001001100;
	ram[110] = 58'b1110011100101010111000011000010011010111000110000111100010;
	ram[111] = 58'b1110011011110110101111011011000000000100111000011101100100;
	ram[112] = 58'b1110011011000010101100010101101101110110100101000001000000;
	ram[113] = 58'b1110011010001110101111000111011011011100110100001011101111;
	ram[114] = 58'b1110011001011010110111101111001001101001111101111110001110;
	ram[115] = 58'b1110011000100111000110001011111001011110100110101011010000;
	ram[116] = 58'b1110010111110011011010011100101101000010110111001010001100;
	ram[117] = 58'b1110010110111111110100100000100100111001111110011001110011;
	ram[118] = 58'b1110010110001100010100010110100010101110101110100000000000;
	ram[119] = 58'b1110010101011000111001111101100111100000100011111000001001;
	ram[120] = 58'b1110010100100101100101010100110111001000101101111100100000;
	ram[121] = 58'b1110010011110010010110011011010011000010010011100110111100;
	ram[122] = 58'b1110010010111111001101001111111101101111100010010111000110;
	ram[123] = 58'b1110010010001100001001110001111001000111001111010101010100;
	ram[124] = 58'b1110010001011001001100000000001001111001001101000110100100;
	ram[125] = 58'b1110010000100110010011111001110001011110011101010111001100;
	ram[126] = 58'b1110001111110011100001011101110011001111110101010011000010;
	ram[127] = 58'b1110001111000000110100101011010011101100100000110010110001;
	ram[128] = 58'b1110001110001110001101100001010110101000000011111000000000;
	ram[129] = 58'b1110001101011011101011111110111111001010100110100001100111;
	ram[130] = 58'b1110001100101001010000000011010001100010011111101000111000;
	ram[131] = 58'b1110001011110110111001101101010011000100000001101101000000;
	ram[132] = 58'b1110001011000100101000111100000111011111001011110000000000;
	ram[133] = 58'b1110001010010010011101101110110011101001110111010110101100;
	ram[134] = 58'b1110001001100000011000000100011101011111100101010111001010;
	ram[135] = 58'b1110001000101110010111111100001000011111001011010010100001;
	ram[136] = 58'b1110000111111100011101010100111011110110100111011111100000;
	ram[137] = 58'b1110000111001010101000001101111011011110110010100101110000;
	ram[138] = 58'b1110000110011000111000100110001110111111001110000000110110;
	ram[139] = 58'b1110000101100111001110011100111010101010100111001100111101;
	ram[140] = 58'b1110000100110101101001110001000101101001100100001011010100;
	ram[141] = 58'b1110000100000100001010100001110110011000111100111000000011;
	ram[142] = 58'b1110000011010010110000101110010011100010010001000110000010;
	ram[143] = 58'b1110000010100001011100010101100011000011011110001010100100;
	ram[144] = 58'b1110000001110000001101010110101100110111010110100111110000;
	ram[145] = 58'b1110000000111111000011110000110111010100111100100100011111;
	ram[146] = 58'b1110000000001101111111100011001010101111110100010011011110;
	ram[147] = 58'b1101111111011101000000101100101101110111110110111111110100;
	ram[148] = 58'b1101111110101100000111001100101001011001001101001100101100;
	ram[149] = 58'b1101111101111011010011000010000100011100011001101100001011;
	ram[150] = 58'b1101111101001010100100001100000111001110001010000000000000;
	ram[151] = 58'b1101111100011001111010101001111010111111000011101110000001;
	ram[152] = 58'b1101111011101001010110011010100110100100100011100110100000;
	ram[153] = 58'b1101111010111000110111011101010100011111000011110010111111;
	ram[154] = 58'b1101111010001000011101110001001100110011110101000100100110;
	ram[155] = 58'b1101111001011000001001010101011000101011110011001101110100;
	ram[156] = 58'b1101111000100111111010001001000000100100010011101110100100;
	ram[157] = 58'b1101110111110111110000001011001111101101000011001011101100;
	ram[158] = 58'b1101110111000111101011011011001110000011100011000000100010;
	ram[159] = 58'b1101110110010111101011111000000110010111011111011111101001;
	ram[160] = 58'b1101110101100111110001100001000010101100110001110110000000;
	ram[161] = 58'b1101110100110111111100010101001101010010111100010001110000;
	ram[162] = 58'b1101110100001000001100010011101111101101111001100001111000;
	ram[163] = 58'b1101110011011000100001011011110101011011101000001111000101;
	ram[164] = 58'b1101110010101000111011101100101000010111001011110000000000;
	ram[165] = 58'b1101110001111001011011000101010100010101011001001011000000;
	ram[166] = 58'b1101110001001001111111100101000011101000010000000010100000;
	ram[167] = 58'b1101110000011010101001001011000010011011001111100110110001;
	ram[168] = 58'b1101101111101011010111110110011010100000001011101011011000;
	ram[169] = 58'b1101101110111100001011100110011010000110111100000001001111;
	ram[170] = 58'b1101101110001101000100011010001010100000111111011000000000;
	ram[171] = 58'b1101101101011110000010010000111000100110101101101111110101;
	ram[172] = 58'b1101101100101111000101001001110001011011011011001000010100;
	ram[173] = 58'b1101101100000000001101000100000000011111111001110100110011;
	ram[174] = 58'b1101101011010001011001111110110001100000001001101011001000;
	ram[175] = 58'b1101101010100010101011111001010010110111001010010000000000;
	ram[176] = 58'b1101101001110100000010110010101111110000001110001011010000;
	ram[177] = 58'b1101101001000101011110101010010110111011111101111111001111;
	ram[178] = 58'b1101101000010110111111011111010011111011100110011111100000;
	ram[179] = 58'b1101100111101000100101010000110100111110110001101010010101;
	ram[180] = 58'b1101100110111010001111111110000111101001010101001100110000;
	ram[181] = 58'b1101100110001011111111100110011000110011011110010111001100;
	ram[182] = 58'b1101100101011101110100001000110111001100110110000001101000;
	ram[183] = 58'b1101100100101111101101100100110000000011000001000100000001;
	ram[184] = 58'b1101100100000001101011111001010010011010101111001000000000;
	ram[185] = 58'b1101100011010011101111000101101100101100111011111011100111;
	ram[186] = 58'b1101100010100101110111001001001100100110111010110001100110;
	ram[187] = 58'b1101100001111000000100000011000000110110101011100111110100;
	ram[188] = 58'b1101100001001010010101110010011001001010101001110000000100;
	ram[189] = 58'b1101100000011100101100010110100011101111011110001001101011;
	ram[190] = 58'b1101011111101111000111101110101111110010001101100000001000;
	ram[191] = 58'b1101011111000001100111111010001100101010001101110110010000;
	ram[192] = 58'b1101011110010100001100111000001001111001000011111101000000;
	ram[193] = 58'b1101011101100110110110100111111000000000010100011111011100;
	ram[194] = 58'b1101011100111001100101001000100101001010001111100100101110;
	ram[195] = 58'b1101011100001100011000011001100011000010011010110101010000;
	ram[196] = 58'b1101011011011111010000011010000000000111011100011100011100;
	ram[197] = 58'b1101011010110010001101001001001110011000110100010101001100;
	ram[198] = 58'b1101011010000101001110100110011100101001010100010001011010;
	ram[199] = 58'b1101011001011000010100110000111100010110101001000100110001;
	ram[200] = 58'b1101011000101011011111100111111110010010101110000000000000;
	ram[201] = 58'b1101010111111110101111001010110010100011111000001001000111;
	ram[202] = 58'b1101010111010010000011011000101011111010101011011011011000;
	ram[203] = 58'b1101010110100101011100010000111001000110010001011000010100;
	ram[204] = 58'b1101010101111000111001110010101110000000000001000111010000;
	ram[205] = 58'b1101010101001100011011111101011010100000000011000000000000;
	ram[206] = 58'b1101010100100000000010110000010000010010111110100100100000;
	ram[207] = 58'b1101010011110011101110001010100010000100001111011110001001;
	ram[208] = 58'b1101010011000111011110001011100000111110011000001100000000;
	ram[209] = 58'b1101010010011011010010110010011111111111110111000000000000;
	ram[210] = 58'b1101010001101111001011111110110000100110010111000000111000;
	ram[211] = 58'b1101010001000011001001101111100101001110001101101111110100;
	ram[212] = 58'b1101010000010111001100000100010000011101001100000000000000;
	ram[213] = 58'b1101001111101011010010111100000101110111010111101001110011;
	ram[214] = 58'b1101001110111111011110010110010111100000001111100010100000;
	ram[215] = 58'b1101001110010011101110010010010111100100110001110110010000;
	ram[216] = 58'b1101001101101000000010101111011010111001110100011100101000;
	ram[217] = 58'b1101001100111100011011101100110011111110110011101011110000;
	ram[218] = 58'b1101001100010000111001001001110110010001010010000101110110;
	ram[219] = 58'b1101001011100101011011000101110100100011010001001100011101;
	ram[220] = 58'b1101001010111010000001100000000100001110000000011010010000;
	ram[221] = 58'b1101001010001110101100010111110111100001000110010001001100;
	ram[222] = 58'b1101001001100011011011101100100100000111110000110100000010;
	ram[223] = 58'b1101001000111000001111011101011011101111010101100100000000;
	ram[224] = 58'b1101001000001101000111101001110101001001011110000010000000;
	ram[225] = 58'b1101000111100010000100010001000011001010000110101101100111;
	ram[226] = 58'b1101000110110111000101010010011011001011100110011101111000;
	ram[227] = 58'b1101000110001100001010101101010001111100101011001010011101;
	ram[228] = 58'b1101000101100001010100100000111011100000100101001110011100;
	ram[229] = 58'b1101000100110110100010101100101100110111110011111110101100;
	ram[230] = 58'b1101000100001011110101001111111011111111110101111110001010;
	ram[231] = 58'b1101000011100001001100001001111101010110010111011010101001;
	ram[232] = 58'b1101000010110110100111011010000111001010001101100100011000;
	ram[233] = 58'b1101000010001100000110111111101110001010100001010010111100;
	ram[234] = 58'b1101000001100001101010111010001000000011010010000001011000;
	ram[235] = 58'b1101000000110111010011001000101011011101000110001101000000;
	ram[236] = 58'b1101000000001100111111101010101100101101000011001001010000;
	ram[237] = 58'b1100111111100010110000011111100011100000110011011100001100;
	ram[238] = 58'b1100111110111000100101100110100101010010100001010110000010;
	ram[239] = 58'b1100111110001110011110111111001000011000110101100101000001;
	ram[240] = 58'b1100111101100100011100101000100011010010110100010000000000;
	ram[241] = 58'b1100111100111010011110100010001101011011101011110010111111;
	ram[242] = 58'b1100111100010000100100101011011011111011101100000001111000;
	ram[243] = 58'b1100111011100110101111000011100110011110110010000111010000;
	ram[244] = 58'b1100111010111100111101101010000011010001110001011000110000;
	ram[245] = 58'b1100111010010011010000011110001011000100101100001001101100;
	ram[246] = 58'b1100111001101001100111011111010011100001001110100011101000;
	ram[247] = 58'b1100111001000000000010101100110101100111101100001100010000;
	ram[248] = 58'b1100111000010110100010000110000111010010010010111000100000;
	ram[249] = 58'b1100110111101101000101101010100000001010100110011111000000;
	ram[250] = 58'b1100110111000011101101011001011000110101101010110001000110;
	ram[251] = 58'b1100110110011010011001010010001001001101000110111001110101;
	ram[252] = 58'b1100110101110001001001010100001001010010100100010000000000;
	ram[253] = 58'b1100110101000111111101011110110000011100011010111000110011;
	ram[254] = 58'b1100110100011110110101110001010110111100011011000010001000;
	ram[255] = 58'b1100110011110101110010001011010101111111011101111010010000;
	ram[256] = 58'b1100110011001100110010101100000101010011111000110000000000;
	ram[257] = 58'b1100110010100011110111010010111110010110010010101100011111;
	ram[258] = 58'b1100110001111010111111111111011001000100110101000111100000;
	ram[259] = 58'b1100110001010010001100110000101110011000101010101101001101;
	ram[260] = 58'b1100110000101001011101100110010111010010110000100111110000;
	ram[261] = 58'b1100110000000000110010011111101101101110110010010111101100;
	ram[262] = 58'b1100101111011000001011011100001010001010001010000010101000;
	ram[263] = 58'b1100101110101111101000011011000101111101000001001110000100;
	ram[264] = 58'b1100101110000111001001011011111010100111001100010111100000;
	ram[265] = 58'b1100101101011110101110011110000001110000001000111100011100;
	ram[266] = 58'b1100101100110110010111100000110101000110111011100010011000;
	ram[267] = 58'b1100101100001110000100100011101110100010001101111110110100;
	ram[268] = 58'b1100101011100101110101100110001000000000001101011111010000;
	ram[269] = 58'b1100101010111101101010100111011011100110101000110001001100;
	ram[270] = 58'b1100101010010101100011100111000011100010101110001010001000;
	ram[271] = 58'b1100101001101101100000100100011010001001001001101111100100;
	ram[272] = 58'b1100101001000101100001011110111001110110000011011111000000;
	ram[273] = 58'b1100101000011101100110010101111100011010011110010110000111;
	ram[274] = 58'b1100100111110101101111001000111101010011111000111110000000;
	ram[275] = 58'b1100100111001101111011110111010111010100100100010000110101;
	ram[276] = 58'b1100100110100110001100100000100100100011101101111101001100;
	ram[277] = 58'b1100100101111110100001000100000000110100101011001111011011;
	ram[278] = 58'b1100100101010110111001100001000111001111100101100101101010;
	ram[279] = 58'b1100100100101111010101110111010010010001100101010101000100;
	ram[280] = 58'b1100100100000111110110000101111110000011100110000000101000;
	ram[281] = 58'b1100100011100000011010001100100101010001001110010000001111;
	ram[282] = 58'b1100100010111001000010001010100011011111100001010010011000;
	ram[283] = 58'b1100100010010001101101111111010101001100110001010100010101;
	ram[284] = 58'b1100100001101010011101101010010110001100001001000000000000;
	ram[285] = 58'b1100100001000011010001001011000000110011110100010111001011;
	ram[286] = 58'b1100100000011100001000100000110010101001010011000011001000;
	ram[287] = 58'b1100011111110101000011101011000111110100111000110011000001;
	ram[288] = 58'b1100011111001110000010101001011011000010000100001110000000;
	ram[289] = 58'b1100011110100111000101011011001010001011000100111110000111;
	ram[290] = 58'b1100011110000000001011111111110000111011010010111101111110;
	ram[291] = 58'b1100011101011001010110010110101011110110111101011101000000;
	ram[292] = 58'b1100011100110010100100011111010111101001001100011100000000;
	ram[293] = 58'b1100011100001011110110011001010001000011111111000011101011;
	ram[294] = 58'b1100011011100101001100000011110101000000001001111011001010;
	ram[295] = 58'b1100011010111110100101011110100000011101010101011110100100;
	ram[296] = 58'b1100011010011000000010101000110000100001111100010101100000;
	ram[297] = 58'b1100011001110001100011100010000010011011001001101001100111;
	ram[298] = 58'b1100011001001011001000001001110011011100110111011101000110;
	ram[299] = 58'b1100011000100100110000011111100001000001101101000001010000;
	ram[300] = 58'b1100010111111110011100100010101000101010111101001101000000;
	ram[301] = 58'b1100010111011000001100010010100111001111001010000100101100;
	ram[302] = 58'b1100010110110001111111101110111011001110011000101100010010;
	ram[303] = 58'b1100010110001011110110110111000010011101110101010100111001;
	ram[304] = 58'b1100010101100101110001101010011010000111111101011001010000;
	ram[305] = 58'b1100010100111111110000001000100001110001110000011100011111;
	ram[306] = 58'b1100010100011001110010010000110101010000010000101101111000;
	ram[307] = 58'b1100010011110011111000000010110101000110101010110011100101;
	ram[308] = 58'b1100010011001110000001011101111110001000011001000100110000;
	ram[309] = 58'b1100010010101000001110100001101110110001110110101001100011;
	ram[310] = 58'b1100010010000010011111001101100110010111000000010000101010;
	ram[311] = 58'b1100010001011100110011100001000011100001000000000000000000;
	ram[312] = 58'b1100010000110111001011011011100100001110010111101001001000;
	ram[313] = 58'b1100010000010001100110111100100111010101001000011101110000;
	ram[314] = 58'b1100001111101100000110000011101011110001101001001001000110;
	ram[315] = 58'b1100001111000110101000110000010001010111011110111100100101;
	ram[316] = 58'b1100001110100001001111000001110111001111100000100000010000;
	ram[317] = 58'b1100001101111011111000110111111011000111001011000000000000;
	ram[318] = 58'b1100001101010110100110010001111101110101101010000011010010;
	ram[319] = 58'b1100001100110001010111001111011110000101110010110001000000;
	ram[320] = 58'b1100001100001100001011101111111011011001011110101011000000;
	ram[321] = 58'b1100001011100111000011110010110101011000110010011111000000;
	ram[322] = 58'b1100001011000001111111010111101011110001111100101010101110;
	ram[323] = 58'b1100001010011100111110011101111111001001111011101110111101;
	ram[324] = 58'b1100001001111000000001000101001101111001111011110111110000;
	ram[325] = 58'b1100001001010011000111001100111001100011101101000000101100;
	ram[326] = 58'b1100001000101110010000110100100000101100101110000100111010;
	ram[327] = 58'b1100001000001001011101111011100101000010101100001011010001;
	ram[328] = 58'b1100000111100100101110100001100101010111010011001110000000;
	ram[329] = 58'b1100000111000000000010100110000010110011101110000101011111;
	ram[330] = 58'b1100000110011011011010001000011101110110100101100000000000;
	ram[331] = 58'b1100000101110110110101001000010111000100011111000000111101;
	ram[332] = 58'b1100000101010010010011100101001111000111111011100101000000;
	ram[333] = 58'b1100000100101101110101011110100110000001000101101001001100;
	ram[334] = 58'b1100000100001001011010110011111101010110100110000011001000;
	ram[335] = 58'b1100000011100101000011100100110110000100100111111001000000;
	ram[336] = 58'b1100000011000000101111110000110001001101001100000000000000;
	ram[337] = 58'b1100000010011100011111010111001111001000000000001101010111;
	ram[338] = 58'b1100000001111000010010010111110001110010111001001110000000;
	ram[339] = 58'b1100000001010100001000110001111001110001001110010101000000;
	ram[340] = 58'b1100000000110000000010100101001001001100010010000000110000;
	ram[341] = 58'b1100000000001011111111110001000001100010111110001010101100;
	ram[342] = 58'b1011111111101000000000010101000011101001111110001001011010;
	ram[343] = 58'b1011111111000100000100010000110001001011101100110011101001;
	ram[344] = 58'b1011111110100000001011100011101100101000000111111001101000;
	ram[345] = 58'b1011111101111100010110001101010111110100111000001111010111;
	ram[346] = 58'b1011111101011000100100001101010011001101101000110101110110;
	ram[347] = 58'b1011111100110100110101100011000010010011000001100010100101;
	ram[348] = 58'b1011111100010001001010001110000111001011100000101100000100;
	ram[349] = 58'b1011111011101101100010001110000010100011110000000100100011;
	ram[350] = 58'b1011111011001001111101100010011000001100110111101110010010;
	ram[351] = 58'b1011111010100110011100001010101001101110010111011111100100;
	ram[352] = 58'b1011111010000010111110000110011010010100100100100110100000;
	ram[353] = 58'b1011111001011111100011010101001011000010011111110000000000;
	ram[354] = 58'b1011111000111100001011110110011111111110111111000111111110;
	ram[355] = 58'b1011111000011000110111101001111010011000000111000101110100;
	ram[356] = 58'b1011110111110101100110101110111110011111011101101010011100;
	ram[357] = 58'b1011110111010010011001000101001110011101100000100101111011;
	ram[358] = 58'b1011110110101111001110101100001101001111101000010011101000;
	ram[359] = 58'b1011110110001100000111100011011101111000100101000001000000;
	ram[360] = 58'b1011110101101001000011101010100011100000011101011110011000;
	ram[361] = 58'b1011110101000110000011000001000001010100101101101111101111;
	ram[362] = 58'b1011110100100011000101100110011010101000000101111101100000;
	ram[363] = 58'b1011110100000000001011011010010010000011011011011000010101;
	ram[364] = 58'b1011110011011101010100011100001100100010100000011101000000;
	ram[365] = 58'b1011110010111010100000101011101100001001100000101101101011;
	ram[366] = 58'b1011110010010111110000001000010101001111011110010001110010;
	ram[367] = 58'b1011110001110101000010110001101011100001011011100001000000;
	ram[368] = 58'b1011110001010010011000100111010010110001100111100001000000;
	ram[369] = 58'b1011110000101111110001101000101110110111011100110110001111;
	ram[370] = 58'b1011110000001101001101110101100011000000100010001110000000;
	ram[371] = 58'b1011101111101010101101001101010011001110101100010011000101;
	ram[372] = 58'b1011101111001000001111101111100101000110101100111011000000;
	ram[373] = 58'b1011101110100101110101011011111011010110101010010110111011;
	ram[374] = 58'b1011101110000011011110010001111010111110100100001110011010;
	ram[375] = 58'b1011101101100001001010010001000111100101101110010101011001;
	ram[376] = 58'b1011101100111110111001011001000110010110001011110010000000;
	ram[377] = 58'b1011101100011100101011101001011011000001011010010101101111;
	ram[378] = 58'b1011101011111010100001000001101010111011011100001001100110;
	ram[379] = 58'b1011101011011000011001100001011001111111110100010011000101;
	ram[380] = 58'b1011101010110110010101001000001100111101110110001000100100;
	ram[381] = 58'b1011101010010100010011110101101010000111000001010100101011;
	ram[382] = 58'b1011101001110010010101101001010100001000100111110100001000;
	ram[383] = 58'b1011101001010000011010100010110001011101111110110000010000;
	ram[384] = 58'b1011101000101110100010100001100110011011100010101000000000;
	ram[385] = 58'b1011101000001100101101100101011000001001010000000001110000;
	ram[386] = 58'b1011100111101010111011101101101100100010011000001110101110;
	ram[387] = 58'b1011100111001001001100111010001000001010000110001001110100;
	ram[388] = 58'b1011100110100111100001001010010000010110111011011010011100;
	ram[389] = 58'b1011100110000101111000011101101010100100001110010011000000;
	ram[390] = 58'b1011100101100100010010110011111101000000011100111010000000;
	ram[391] = 58'b1011100101000010110000001100101011110011111001101001000001;
	ram[392] = 58'b1011100100100001010000100111011110000100111000101010111000;
	ram[393] = 58'b1011100011111111110100000011111000110011100100011010110111;
	ram[394] = 58'b1011100011011110011010100001100001110011001010110101110110;
	ram[395] = 58'b1011100010111101000011111111111110001101011110011100110100;
	ram[396] = 58'b1011100010011011110000011110110101011011011110001111010000;
	ram[397] = 58'b1011100001111010011111111101101100110000010011111110101100;
	ram[398] = 58'b1011100001011001010010011100001010010010000000011010001000;
	ram[399] = 58'b1011100000111000000111111001110100001011001110010100000100;
	ram[400] = 58'b1011100000010111000000010110010000101011010001011111000000;
	ram[401] = 58'b1011011111110101111011110001000101011000001000011110000111;
	ram[402] = 58'b1011011111010100111010001001111010000110010010101100011110;
	ram[403] = 58'b1011011110110011111011100000010011110111000000001101000000;
	ram[404] = 58'b1011011110010010111111110011111001111001111011110011101100;
	ram[405] = 58'b1011011101110010000111000100010010110101010110111011101100;
	ram[406] = 58'b1011011101010001010001010001000101010100000101101111101010;
	ram[407] = 58'b1011011100110000011110011001110111010111101101010100000001;
	ram[408] = 58'b1011011100001111101110011110010000100001111001100001101000;
	ram[409] = 58'b1011011011101111000001011101110111101011000001000101111111;
	ram[410] = 58'b1011011011001110010111011000010011101111111001010100100110;
	ram[411] = 58'b1011011010101101110000001101001011000100001100110000110100;
	ram[412] = 58'b1011011010001101001011111100000100101101110001011010010000;
	ram[413] = 58'b1011011001101100101010100100101001010010000010111011000011;
	ram[414] = 58'b1011011001001100001100000110011110100100011100001110010010;
	ram[415] = 58'b1011011000101011110000100001001011111000000100000011000100;
	ram[416] = 58'b1011011000001011010111110100011001010001111000011101100000;
	ram[417] = 58'b1011010111101011000001111111101110001101101010101011110000;
	ram[418] = 58'b1011010111001010101111000010110000110000101101110011001110;
	ram[419] = 58'b1011010110101010011110111101001010100111110101111010000101;
	ram[420] = 58'b1011010110001010010001101110100010000001000010101111000000;
	ram[421] = 58'b1011010101101010000111010110011110101001100001101100000000;
	ram[422] = 58'b1011010101001001111111110100101000010010110010111001111010;
	ram[423] = 58'b1011010100101001111011001000100111011111111001100001000100;
	ram[424] = 58'b1011010100001001111001010010000011011101100100011000000000;
	ram[425] = 58'b1011010011101001111010010000100100110111010100001010011100;
	ram[426] = 58'b1011010011001001111110000011110011000010011011001001110110;
	ram[427] = 58'b1011010010101010000100101011010110000101101010111100000101;
	ram[428] = 58'b1011010010001010001110000110110110001100000010011001010000;
	ram[429] = 58'b1011010001101010011010010101111100010001110001101101000011;
	ram[430] = 58'b1011010001001010101001011000001111111101000111000111000010;
	ram[431] = 58'b1011010000101010111011001101011000111000100011101101100001;
	ram[432] = 58'b1011010000001011001111110101000001100110110101000000000000;
	ram[433] = 58'b1011001111101011100111001110110000100000101101001011100111;
	ram[434] = 58'b1011001111001100000001011010001110110111001001000101001110;
	ram[435] = 58'b1011001110101100011110010111000101010010001011110111010100;
	ram[436] = 58'b1011001110001100111110000100111101001010110101110001001100;
	ram[437] = 58'b1011001101101101100000100011011101110111100101110001101100;
	ram[438] = 58'b1011001101001110000101110010010000111001100111011010000000;
	ram[439] = 58'b1011001100101110101101110000111111110110000010001111100100;
	ram[440] = 58'b1011001100001111011000011111010010001111101011000100100000;
	ram[441] = 58'b1011001011110000000101111100110010100000011100011111111100;
	ram[442] = 58'b1011001011010000110110001001001000010011010110000000000000;
	ram[443] = 58'b1011001010110001101001000011111101011101100001101111100101;
	ram[444] = 58'b1011001010010010011110101100111011001011011010000111100100;
	ram[445] = 58'b1011001001110011010111000011101010101101010111101010110000;
	ram[446] = 58'b1011001001010100010010000111110100101011001100111101110010;
	ram[447] = 58'b1011001000110101001111111001000011110110010101000000000100;
	ram[448] = 58'b1011001000010110010000010111000000010001111000111001000000;
	ram[449] = 58'b1011000111110111010011100001010100001010100100101011100111;
	ram[450] = 58'b1011000111011000011001010111101001000100011010111110000000;
	ram[451] = 58'b1011000110111001100001111001100111111010111101101011111101;
	ram[452] = 58'b1011000110011010101101000110111011110010110101111111110000;
	ram[453] = 58'b1011000101111011111010111111001100010110100111111100101100;
	ram[454] = 58'b1011000101011101001011100010000101011110111100011110101000;
	ram[455] = 58'b1011000100111110011110101111001111101010100001010001000000;
	ram[456] = 58'b1011000100011111110100100110010101100000111000011101111000;
	ram[457] = 58'b1011000100000001001101000111000000010100110100010111110000;
	ram[458] = 58'b1011000011100010101000010000111010110101011010011111011000;
	ram[459] = 58'b1011000011000100000110000011101110011101000110011011110100;
	ram[460] = 58'b1011000010100101100110011111000110000010011110000100110100;
	ram[461] = 58'b1011000010000111001001100010101011110011101001101110101011;
	ram[462] = 58'b1011000001101000101111001110001001010110011100111111110010;
	ram[463] = 58'b1011000001001010010111100001001001000000100101000110101001;
	ram[464] = 58'b1011000000101100000010011011010101110111011110011011000000;
	ram[465] = 58'b1011000000001101101111111100011001101100001101010011101111;
	ram[466] = 58'b1010111111101111100000000011111111101011100100110001001110;
	ram[467] = 58'b1010111111010001010010110001110001101110000101100110111101;
	ram[468] = 58'b1010111110110011001000000101011010011011111100101110101100;
	ram[469] = 58'b1010111110010100111111111110100101001100111001000011001100;
	ram[470] = 58'b1010111101110110111010011100111100000100100000000110011010;
	ram[471] = 58'b1010111101011000110111100000001010100001101111010001101001;
	ram[472] = 58'b1010111100111010110111000111111010000011101111010010100000;
	ram[473] = 58'b1010111100011100111001010011110110111100011110011100000000;
	ram[474] = 58'b1010111011111110111110000011101011011110001000100110000000;
	ram[475] = 58'b1010111011100001000101010111000010101010010010111011110100;
	ram[476] = 58'b1010111011000011001111001101101000010001110010001001100100;
	ram[477] = 58'b1010111010100101011011100111000110110001100110010011001100;
	ram[478] = 58'b1010111010000111101010100011001000101010011010110000001000;
	ram[479] = 58'b1010111001101001111100000001011010100011010011000010010001;
	ram[480] = 58'b1010111001001100010000000001100111000011111101000010000000;
	ram[481] = 58'b1010111000101110100110100011011010001110110001011010111100;
	ram[482] = 58'b1010111000010000111111100110011110000111000100010001111110;
	ram[483] = 58'b1010110111110011011011001010011110110110010000000111010100;
	ram[484] = 58'b1010110111010101111001001111000111111101101011100001011100;
	ram[485] = 58'b1010110110111000011001110100000101101101100101000111111011;
	ram[486] = 58'b1010110110011010111100111001000010010111011010000000000000;
	ram[487] = 58'b1010110101111101100010011101101010010010010100100110110001;
	ram[488] = 58'b1010110101100000001010100001101001001101100000000000000000;
	ram[489] = 58'b1010110101000010110101000100101011100110110100111100000000;
	ram[490] = 58'b1010110100100101100010000110011011111101101101101101110110;
	ram[491] = 58'b1010110100001000010001100110100110110110111001001011010000;
	ram[492] = 58'b1010110011101011000011100100110111100011111110010100000000;
	ram[493] = 58'b1010110011001101111000000000111011011011100100111100110011;
	ram[494] = 58'b1010110010110000101110111010011101110110000010001000000000;
	ram[495] = 58'b1010110010010011101000010001001010001111001001100011100100;
	ram[496] = 58'b1010110001110110100100000100101101011100010111010001000000;
	ram[497] = 58'b1010110001011001100010010100110011101011010010000001110000;
	ram[498] = 58'b1010110000111100100011000001001001001100110101010111100000;
	ram[499] = 58'b1010110000011111100110001001011001101010010001000110000101;
	ram[500] = 58'b1010110000000010101011101101010010000110001100000000000000;
	ram[501] = 58'b1010101111100101110011101100011110111011011100001001010011;
	ram[502] = 58'b1010101111001000111110000110101011111101001110111000011010;
	ram[503] = 58'b1010101110101100001010111011100110010111111100000011000001;
	ram[504] = 58'b1010101110001111011010001010111010110000001101111101001000;
	ram[505] = 58'b1010101101110010101011110100010101101101111110101010010111;
	ram[506] = 58'b1010101101010101111111110111100011010001100100010110011000;
	ram[507] = 58'b1010101100111001010110010100010000001001011100101011010000;
	ram[508] = 58'b1010101100011100101111001010001001110010000011001001000000;
	ram[509] = 58'b1010101100000000001010011000111101000000001011011111101100;
	ram[510] = 58'b1010101011100011101000000000010110000001001001011110000010;
	ram[511] = 58'b1010101011000111001000000000000010011010111001011010100100;
	ram[512] = 58'b1010101010101010101010010111101110100001001010000000000000;
	ram[513] = 58'b1010101010001110001111000111001000000000001001111101110000;
	ram[514] = 58'b1010101001110001110110001101111011010010000000010000101110;
	ram[515] = 58'b1010101001010101011111101011110110001001001011010101000000;
	ram[516] = 58'b1010101000111001001011100000100101000110000111110111000000;
	ram[517] = 58'b1010101000011100111001101011110101010111000001100011101011;
	ram[518] = 58'b1010101000000000101010001101010100110111101001101000000000;
	ram[519] = 58'b1010100111100100011101000100110000010001111000010000000000;
	ram[520] = 58'b1010100111001000010010010001110100111101001101010001111000;
	ram[521] = 58'b1010100110101100001001110100010000111110100111010001110000;
	ram[522] = 58'b1010100110010000000011101011110001001001010011110110000000;
	ram[523] = 58'b1010100101110011111111111000000011101000010110111111010100;
	ram[524] = 58'b1010100101010111111110011000110100101010110101111101000000;
	ram[525] = 58'b1010100100111011111111001101110011001100001110111100110000;
	ram[526] = 58'b1010100100100000000010010110101100001100000011100111100010;
	ram[527] = 58'b1010100100000100000111110011001110000001011011100100000000;
	ram[528] = 58'b1010100011101000001111100011000101000111110001101101110000;
	ram[529] = 58'b1010100011001100011001100110000000100110011100000000000000;
	ram[530] = 58'b1010100010110000100101111011101101101001000101111011111000;
	ram[531] = 58'b1010100010010100110100100011111010001000101000111100000101;
	ram[532] = 58'b1010100001111001000101011110010100000000111100111101001100;
	ram[533] = 58'b1010100001011101011000101010101001111010111100001010001011;
	ram[534] = 58'b1010100001000001101110001000101000100100001111110010001010;
	ram[535] = 58'b1010100000100110000101110111111111010101101110010101010001;
	ram[536] = 58'b1010100000001010011111111000011011000011000001000101101000;
	ram[537] = 58'b1010011111101110111100001001101011001010101111010001000111;
	ram[538] = 58'b1010011111010011011010101011011100100110011111011001010110;
	ram[539] = 58'b1010011110110111111011011101011110111010100111010110111101;
	ram[540] = 58'b1010011110011100011110011111011111110000100000100000010000;
	ram[541] = 58'b1010011110000001000011110001001100110100100100100110100011;
	ram[542] = 58'b1010011101100101101011010010010101110011101010011110001000;
	ram[543] = 58'b1010011101001010010101000010100111110110000111100111001001;
	ram[544] = 58'b1010011100101111000001000001110010101110011011011110000000;
	ram[545] = 58'b1010011100010011101111001111100011101010110000101000011111;
	ram[546] = 58'b1010011011111000011111101011101001111001011110110100101110;
	ram[547] = 58'b1010011011011101010010010101110100000010000000101001010000;
	ram[548] = 58'b1010011011000010000111001101110000101110100101101111000000;
	ram[549] = 58'b1010011010100110111110010011001110101100010010001011010011;
	ram[550] = 58'b1010011010001011110111100101111100000001010110111000101000;
	ram[551] = 58'b1010011001110000110011000101101000110011101111010000101001;
	ram[552] = 58'b1010011001010101110000110010000010100101101100110110000000;
	ram[553] = 58'b1010011000111010110000101010111000111001000111000111000000;
	ram[554] = 58'b1010011000011111110010101111111010101001000000000010100110;
	ram[555] = 58'b1010011000000100110111000000110110001001101100010010110100;
	ram[556] = 58'b1010010111101001111101011101011011000101010001010100000000;
	ram[557] = 58'b1010010111001111000110000101011000011111000010110010110011;
	ram[558] = 58'b1010010110110100010000111000011101011101000011101001010010;
	ram[559] = 58'b1010010110011001011101110110011000011110101110000011100001;
	ram[560] = 58'b1010010101111110101100111110111001011000111101010000000000;
	ram[561] = 58'b1010010101100011111110010001101110110000101010110010001111;
	ram[562] = 58'b1010010101001001010001101110101000100000001001100011111110;
	ram[563] = 58'b1010010100101110100111010101010101111011000001011111110100;
	ram[564] = 58'b1010010100010011111111000101100101101110010110111001001100;
	ram[565] = 58'b1010010011111001011000111111000111111100011100001111100011;
	ram[566] = 58'b1010010011011110110101000001101100000000111011111110101000;
	ram[567] = 58'b1010010011000100010011001101000000000111110110000111100100;
	ram[568] = 58'b1010010010101001110011100000110101101101101110100010000000;
	ram[569] = 58'b1010010010001111010101111100111011000011111001111010011100;
	ram[570] = 58'b1010010001110100111010100000111111110000101110100110000000;
	ram[571] = 58'b1010010001011010100001001100110100000110001111011110010101;
	ram[572] = 58'b1010010001000000001010000000000111101111111110000111000100;
	ram[573] = 58'b1010010000100101110100111010101001110011000010100010100011;
	ram[574] = 58'b1010010000001011100001111100001010000000010001100010100010;
	ram[575] = 58'b1010001111110001010001000100011000110100000011011001000000;
	ram[576] = 58'b1010001111010111000010010011000101011011011000000111000000;
	ram[577] = 58'b1010001110111100110101100111111111101110110101011111111100;
	ram[578] = 58'b1010001110100010101011000010111000010010011110110111100000;
	ram[579] = 58'b1010001110001000100010100011011110011011000111000011110100;
	ram[580] = 58'b1010001101101110011100001001100010110001110110000101111100;
	ram[581] = 58'b1010001101010100010111110100110100110000101000111010110000;
	ram[582] = 58'b1010001100111010010101100101000100011100111000000001011010;
	ram[583] = 58'b1010001100100000010101011010000001111110011101110110000100;
	ram[584] = 58'b1010001100000110010111010011011110001000100101100111100000;
	ram[585] = 58'b1010001011101100011011010001001000011111011010011110111100;
	ram[586] = 58'b1010001011010010100001010010110001010010011010100000011000;
	ram[587] = 58'b1010001010111000101001011000001001011100001101111100101101;
	ram[588] = 58'b1010001010011110110011100000111111111111111101000001110100;
	ram[589] = 58'b1010001010000100111111101101000110100101110111010000110000;
	ram[590] = 58'b1010001001101011001101111100001100111110101110010010010010;
	ram[591] = 58'b1010001001010001011110001110000100001110111111100001110001;
	ram[592] = 58'b1010001000110111110000100010011011100011111010001100000000;
	ram[593] = 58'b1010001000011110000100111001000100000110110111111100101111;
	ram[594] = 58'b1010001000000100011011010001101111000011101001010000101110;
	ram[595] = 58'b1010000111101010110011101100001100010111011001110111100101;
	ram[596] = 58'b1010000111010001001110001000001100000001110111111110110000;
	ram[597] = 58'b1010000110110111101010100101011111111110100001000011000000;
	ram[598] = 58'b1010000110011110001001000011111000010001110111100011101000;
	ram[599] = 58'b1010000110000100101001100011000101101011010101100000010000;
	ram[600] = 58'b1010000101101011001100000010111000111100101110101110100000;
	ram[601] = 58'b1010000101010001110000100011000010111010010000011100000000;
	ram[602] = 58'b1010000100111000010111000011010100011010100000110000011000;
	ram[603] = 58'b1010000100011110111111100011011110010110011110001111010000;
	ram[604] = 58'b1010000100000101101010000011010001101001011111011010010000;
	ram[605] = 58'b1010000011101100010110100010011111010001010010010011000000;
	ram[606] = 58'b1010000011010011000101000000111000001101111011111101001000;
	ram[607] = 58'b1010000010111001110101011110001101100001111000000000010000;
	ram[608] = 58'b1010000010100000100111111010001111101001101111101110100000;
	ram[609] = 58'b1010000010000111011100010100110000111100111101001101011111;
	ram[610] = 58'b1010000001101110010010101101100001111100110010101110001110;
	ram[611] = 58'b1010000001010101001011000100010011001100111110001011110100;
	ram[612] = 58'b1010000000111100000101011000110110100011101011111000011100;
	ram[613] = 58'b1010000000100011000001101010111101010001010101010110110000;
	ram[614] = 58'b1010000000001001111111111010011000101000100111011110011010;
	ram[615] = 58'b1001111111110001000000000110111001111110100001111110000100;
	ram[616] = 58'b1001111111011000000010010000010010000010011011010001100000;
	ram[617] = 58'b1001111110111111000110010110010010110101110110100110111100;
	ram[618] = 58'b1001111110100110001100011000101101110100101010000001011000;
	ram[619] = 58'b1001111110001101010100010111010100011100111100100101110100;
	ram[620] = 58'b1001111101110100011110010001111000001111000101111101010000;
	ram[621] = 58'b1001111101011011101010001000001010000101111010000011011011;
	ram[622] = 58'b1001111101000010110111111001111100001110001000000000000000;
	ram[623] = 58'b1001111100101010000111100111000000001110110111000010011001;
	ram[624] = 58'b1001111100010001011001001111000111001001101110000000010000;
	ram[625] = 58'b1001111011111000101100110010000011010010000100001001001111;
	ram[626] = 58'b1001111011100000000010001111100110010101101100010100101110;
	ram[627] = 58'b1001111011000111011001100111100001011100111100010001010100;
	ram[628] = 58'b1001111010101110110010111001100111000001101111100111101100;
	ram[629] = 58'b1001111010010110001110000101101000010000111001000011000011;
	ram[630] = 58'b1001111001111101101011001011011000010000010000111110100000;
	ram[631] = 58'b1001111001100101001010001010100111000001110111001100000001;
	ram[632] = 58'b1001111001001100101011000011001000010111011101001011001000;
	ram[633] = 58'b1001111000110100001101110100101100111111000100011000011100;
	ram[634] = 58'b1001111000011011110010011111000110111000000101110110000000;
	ram[635] = 58'b1001111000000011011001000010001000101011100011001011110100;
	ram[636] = 58'b1001110111101011000001011101100011110101100111101011100100;
	ram[637] = 58'b1001110111010010101011110001001011000011100101100011000000;
	ram[638] = 58'b1001110110111010010111111100110000011101010111101010010010;
	ram[639] = 58'b1001110110100010000110000000000101100101101000110110110001;
	ram[640] = 58'b1001110110001001110101111010111100101000101001100000000000;
	ram[641] = 58'b1001110101110001100111101101001000011100000111010001001111;
	ram[642] = 58'b1001110101011001011011010110011010101001001000111110011110;
	ram[643] = 58'b1001110101000001010000110110100110001001100111110100000101;
	ram[644] = 58'b1001110100101001001000001101011100101010111011000111000000;
	ram[645] = 58'b1001110100010001000001011010110001001011000101101101010011;
	ram[646] = 58'b1001110011111000111100011110010101011011101110000100001010;
	ram[647] = 58'b1001110011100000111001010111111011110111110010101010010000;
	ram[648] = 58'b1001110011001000111000000111010111100011100001101100111000;
	ram[649] = 58'b1001110010110000111000101100011010010110110101010011100111;
	ram[650] = 58'b1001110010011000111011000110110110110010111001101000011000;
	ram[651] = 58'b1001110010000000111111010110011111011010111110010110110100;
	ram[652] = 58'b1001110001101001000101011011000111011011011100001001010000;
	ram[653] = 58'b1001110001010001001101010100100001011011100100101111101100;
	ram[654] = 58'b1001110000111001010111000010011110110110101000100000100000;
	ram[655] = 58'b1001110000100001100010100100110011100110001000001101100100;
	ram[656] = 58'b1001110000001001101111111011010001110000011101010101110000;
	ram[657] = 58'b1001101111110001111111000101101100000101000110010110101111;
	ram[658] = 58'b1001101111011010010000000011110101111100011110111110001110;
	ram[659] = 58'b1001101111000010100010110101100000111100001101101000000101;
	ram[660] = 58'b1001101110101010110111011010100001000111101001110000001100;
	ram[661] = 58'b1001101110010011001101110010101000101111010111100011000000;
	ram[662] = 58'b1001101101111011100101111101101011010011101101010111111010;
	ram[663] = 58'b1001101101100011111111111011011010100010011100011001000000;
	ram[664] = 58'b1001101101001100011011101011101010100110101101100000101000;
	ram[665] = 58'b1001101100110100111001001110001101010010010101000101110000;
	ram[666] = 58'b1001101100011101011000100010110110110100010010110001110110;
	ram[667] = 58'b1001101100000101111001101001011001101001001011001111101101;
	ram[668] = 58'b1001101011101110011100100001101000110110010011111001000000;
	ram[669] = 58'b1001101011010111000001001011010111100010111111000001001100;
	ram[670] = 58'b1001101010111111100111100110011001011111000110001000000000;
	ram[671] = 58'b1001101010101000001111110010100000101000011101101110010000;
	ram[672] = 58'b1001101010010000111001101111100000110010111000100101100000;
	ram[673] = 58'b1001101001111001100101011101001101110011111111010010111100;
	ram[674] = 58'b1001101001100010010010111011011001101111100001100111101110;
	ram[675] = 58'b1001101001001011000010001001111000011110111111001000110101;
	ram[676] = 58'b1001101000110011110011001000011101111101101100011110111100;
	ram[677] = 58'b1001101000011100100101110110111100010101010000111101011011;
	ram[678] = 58'b1001101000000101011010010101001000001011010100111111111010;
	ram[679] = 58'b1001100111101110010000100010110011101101011001000001000001;
	ram[680] = 58'b1001100111010111001000011111110010111110010101101001100000;
	ram[681] = 58'b1001100111000000000010001011111001011100011100000000000000;
	ram[682] = 58'b1001100110101000111101100110111011001110001110100111011000;
	ram[683] = 58'b1001100110010001111010110000101010101000111010111010110100;
	ram[684] = 58'b1001100101111010111001101000111011110110110100001010010100;
	ram[685] = 58'b1001100101100011111010001111100001110111010101011100001100;
	ram[686] = 58'b1001100101001100111100100100010001011110110000101100000010;
	ram[687] = 58'b1001100100110110000000100110111101110000001100101100110001;
	ram[688] = 58'b1001100100011111000110010111011001110000101100011001010000;
	ram[689] = 58'b1001100100001000001101110101011010011001111011010111010111;
	ram[690] = 58'b1001100011110001010111000000110010001110011000110001111110;
	ram[691] = 58'b1001100011011010100001111001010101100101001000101110110100;
	ram[692] = 58'b1001100011000011101110011110110111101010101001000000001100;
	ram[693] = 58'b1001100010101100111100110001001101011111101101100100110000;
	ram[694] = 58'b1001100010010110001100110000001001101110010011001011101010;
	ram[695] = 58'b1001100001111111011110011011100000110100101001011110001001;
	ram[696] = 58'b1001100001101000110001110011000110101100101000101100100000;
	ram[697] = 58'b1001100001010010000110110110101111010001111100000010111100;
	ram[698] = 58'b1001100000111011011101100110001101111011111111010110000000;
	ram[699] = 58'b1001100000100100110110000001010111010000001000000110001101;
	ram[700] = 58'b1001100000001110010000000111111111001111011000111000000100;
	ram[701] = 58'b1001011111110111101011111001111001010110100111110101101011;
	ram[702] = 58'b1001011111100001001001010110111010110110011000010011110010;
	ram[703] = 58'b1001011111001010101000011110110110000011001011001100010000;
	ram[704] = 58'b1001011110110100001001010001100000110110111101111101000000;
	ram[705] = 58'b1001011110011101101011101110101110001111110011011111000000;
	ram[706] = 58'b1001011110000111001111110110010010111111001111001011100000;
	ram[707] = 58'b1001011101110000110101101000000010101100110011011000010100;
	ram[708] = 58'b1001011101011010011101000011110010001101011111111001111100;
	ram[709] = 58'b1001011101000100000110001001010101110010001011010110011011;
	ram[710] = 58'b1001011100101101110000111000100001000111101001100110001010;
	ram[711] = 58'b1001011100010111011101010001001001001000000010110100100100;
	ram[712] = 58'b1001011100000001001011010011000001100011101010010111111000;
	ram[713] = 58'b1001011011101010111010111101111111011000000001110011010111;
	ram[714] = 58'b1001011011010100101100010001110110111110100110100110000000;
	ram[715] = 58'b1001011010111110011111001110011100001100111000111101100101;
	ram[716] = 58'b1001011010101000010011110011100011011111110100101101000000;
	ram[717] = 58'b1001011010010010001010000001000010100001010001111110000011;
	ram[718] = 58'b1001011001111100000001110110101100000000101010000111100010;
	ram[719] = 58'b1001011001100101111011010100010101101011001011111000010000;
	ram[720] = 58'b1001011001001111110110011001110100000100011111101100000000;
	ram[721] = 58'b1001011000111001110011000110111011001100010110111101011100;
	ram[722] = 58'b1001011000100011110001011011011111101001110100100001111000;
	ram[723] = 58'b1001011000001101110001010111010110101011000101101010111101;
	ram[724] = 58'b1001010111110111110010111010010100111010011110010100001100;
	ram[725] = 58'b1001010111100001110110000100001110011110011111110001000011;
	ram[726] = 58'b1001010111001011111010110100111000000100110110010100001010;
	ram[727] = 58'b1001010110110110000001001100000110011100110111010110100001;
	ram[728] = 58'b1001010110100000001001001001101111100010010011010010101000;
	ram[729] = 58'b1001010110001010010010101101100110010111100011111100011100;
	ram[730] = 58'b1001010101110100011101110111100000111011101001100000011000;
	ram[731] = 58'b1001010101011110101010100111010011011111000100010101000000;
	ram[732] = 58'b1001010101001000111000111100110010111001010101001001000000;
	ram[733] = 58'b1001010100110011001000110111110100101000110110101000110011;
	ram[734] = 58'b1001010100011101011010011000001101000011000100001000000000;
	ram[735] = 58'b1001010100000111101101011101110001101001100100010000000000;
	ram[736] = 58'b1001010011110010000010001000010110110101000011000010000000;
	ram[737] = 58'b1001010011011100011000010111110001100101000101010100111100;
	ram[738] = 58'b1001010011000110110000001011110110111010110110000011100000;
	ram[739] = 58'b1001010010110001001001100100011100011110010000000011000101;
	ram[740] = 58'b1001010010011011100100100001010110101110011101011111000000;
	ram[741] = 58'b1001010010000110000001000010011010110001011010100010011011;
	ram[742] = 58'b1001010001110000011111000111011110010011101110000011101010;
	ram[743] = 58'b1001010001011010111110110000010101010100010001101101100100;
	ram[744] = 58'b1001010001000101011111111100110110000111111001111101100000;
	ram[745] = 58'b1001010000110000000010101100110101010101110000000111110000;
	ram[746] = 58'b1001010000011010100111000000001000001011100111000110000000;
	ram[747] = 58'b1001010000000101001100110110100100011101110100110010111101;
	ram[748] = 58'b1001001111101111110100001111111110111000010001010101000000;
	ram[749] = 58'b1001001111011010011101001100001100001000011101110001101100;
	ram[750] = 58'b1001001111000101000111101011000010101100010100010010110010;
	ram[751] = 58'b1001001110101111110011101100010111111001010011100111001001;
	ram[752] = 58'b1001001110011010100001001111111111111100101100000100000000;
	ram[753] = 58'b1001001110000101010000010101110000110011111111100111000111;
	ram[754] = 58'b1001001101110000000000111101100000011110001100111111101110;
	ram[755] = 58'b1001001101011010110011000111000011110010000101111110100101;
	ram[756] = 58'b1001001101000101100110110010001111101000000011010110110000;
	ram[757] = 58'b1001001100110000011011111110111010101000011000110110101100;
	ram[758] = 58'b1001001100011011010010101100111001101110011111010010100000;
	ram[759] = 58'b1001001100000110001010111100000010011100000100010000000000;
	ram[760] = 58'b1001001011110001000100101100001010010100010101011100100000;
	ram[761] = 58'b1001001011011011111111111101000110111100000000011011111100;
	ram[762] = 58'b1001001011000110111100101110101101111001010010011000000000;
	ram[763] = 58'b1001001010110001111011000000110100110011110111101111010000;
	ram[764] = 58'b1001001010011100111010110011010001111001100100100110000100;
	ram[765] = 58'b1001001010000111111100000101111001101011110001000011110011;
	ram[766] = 58'b1001001001110010111110111000100010011011001111101100110010;
	ram[767] = 58'b1001001001011110000011001011000001110101100111101001110001;
	ram[768] = 58'b1001001001001001001000111101001101101001111110000100000000;
	ram[769] = 58'b1001001000110100010000001110111011101000110101110100010111;
	ram[770] = 58'b1001001000011111011001000000000001100100001111010010011110;
	ram[771] = 58'b1001001000001010100011010000010101001111101000000011110101;
	ram[772] = 58'b1001000111110101101110111111101100011111111010101010111100;
	ram[773] = 58'b1001000111100000111100001101111101001011011110010110011011;
	ram[774] = 58'b1001000111001100001010111010111101001010000110110000001010;
	ram[775] = 58'b1001000110110111011011000110100001110000101001100100000000;
	ram[776] = 58'b1001000110100010101100110000100010000010101000011011100000;
	ram[777] = 58'b1001000110001101111111111000110010110011010111011011100111;
	ram[778] = 58'b1001000101111001010100011111001011001001001010010011110110;
	ram[779] = 58'b1001000101100100101010100011011111111010010000111111110100;
	ram[780] = 58'b1001000101010000000010000101100111101011011100000111010100;
	ram[781] = 58'b1001000100111011011011000101011000011110011111010101001100;
	ram[782] = 58'b1001000100100110110101100010101000010110101000101010110010;
	ram[783] = 58'b1001000100010010010001011101001100110100010000100011110001;
	ram[784] = 58'b1001000011111101101110110100111101000101111010000111000000;
	ram[785] = 58'b1001000011101001001101101001101110001010100010101111000000;
	ram[786] = 58'b1001000011010100101101111011010110101111001111011011100000;
	ram[787] = 58'b1001000011000000001111101001101100111110001110100101010100;
	ram[788] = 58'b1001000010101011110010110100100110011110111110001010001100;
	ram[789] = 58'b1001000010010111010111011011111010100110110010001101010011;
	ram[790] = 58'b1001000010000010111101011111011110011011110001101011101000;
	ram[791] = 58'b1001000001101110100100111111001000110001110110011111011001;
	ram[792] = 58'b1001000001011010001101111010101111010110000101000100101000;
	ram[793] = 58'b1001000001000101111000010010001000111111000100010010110111;
	ram[794] = 58'b1001000000110001100100000101001100000000101100001000110110;
	ram[795] = 58'b1001000000011101010001010011101110110000001011100111001101;
	ram[796] = 58'b1001000000001000111111111101100111100100001000011111100100;
	ram[797] = 58'b1000111111110100110000000010101100010000100001100100110000;
	ram[798] = 58'b1000111111100000100001100010110011110010101010100010110010;
	ram[799] = 58'b1000111111001100010100011101110100000001010001011101111001;
	ram[800] = 58'b1000111110111000001000110011100011111100010011110011100000;
	ram[801] = 58'b1000111110100011111110100011111010000001000111000011001111;
	ram[802] = 58'b1000111110001111110101101110101100101110010101111100111110;
	ram[803] = 58'b1000111101111011101110010011110010000000001010010010110100;
	ram[804] = 58'b1000111101100111101000010011000000111011110010010100011100;
	ram[805] = 58'b1000111101010011100011101100001111100000000100011001001011;
	ram[806] = 58'b1000111100111111100000011111010100110100110101101011011010;
	ram[807] = 58'b1000111100101011011110101100000111011111011001011000110001;
	ram[808] = 58'b1000111100010111011110010010011101100010100110110110000000;
	ram[809] = 58'b1000111100000011011111010010001110001010001011111010001111;
	ram[810] = 58'b1000111011101111100001101011001111011011101010001000010110;
	ram[811] = 58'b1000111011011011100101011101011000100101010100000100010101;
	ram[812] = 58'b1000111011000111101010101000011111101111010100010100000000;
	ram[813] = 58'b1000111010110011110001001100011100001010100001011111111011;
	ram[814] = 58'b1000111010011111111001001001000100100101010111010010000000;
	ram[815] = 58'b1000111010001100000010011110001111001011111100010000000000;
	ram[816] = 58'b1000111001111000001101001011110011010010111010111101000000;
	ram[817] = 58'b1000111001100100011001010001100111001001000001001111001111;
	ram[818] = 58'b1000111001010000100110101111100001100001110111010001101110;
	ram[819] = 58'b1000111000111100110101100101011001110101111001101011011101;
	ram[820] = 58'b1000111000101001000101110011000110111011010000010111101100;
	ram[821] = 58'b1000111000010101010111011000011111000101110100000010110000;
	ram[822] = 58'b1000111000000001101010010101011001110001110001010111011010;
	ram[823] = 58'b1000110111101101111110101001101101010101100101101000111001;
	ram[824] = 58'b1000110111011010010100010101010000101100100000000000000000;
	ram[825] = 58'b1000110111000110101011010111111011010110011011000010000111;
	ram[826] = 58'b1000110110110011000011110001100011101101101000101111110110;
	ram[827] = 58'b1000110110011111011101100010000001010100100001100101001101;
	ram[828] = 58'b1000110110001011111000101001001010100111111001100001000000;
	ram[829] = 58'b1000110101111000010101000110110111001100100101101100100011;
	ram[830] = 58'b1000110101100100110010111010111101100001111011011110110010;
	ram[831] = 58'b1000110101010001010010000101010100101011111000000101100100;
	ram[832] = 58'b1000110100111101110010100101110100010010111010000011000000;
	ram[833] = 58'b1000110100101010010100011100010010111010000111000101001111;
	ram[834] = 58'b1000110100010110110111101000100111101001001000001110000000;
	ram[835] = 58'b1000110100000011011100001010101010001100000011111000100101;
	ram[836] = 58'b1000110011110000000010000010010001001001101101111001111100;
	ram[837] = 58'b1000110011011100101001001111010100010000100110000100101011;
	ram[838] = 58'b1000110011001001010001110001101010001001111110000110100000;
	ram[839] = 58'b1000110010110101111011101001001010000011100100010100000100;
	ram[840] = 58'b1000110010100010100110110101101011001100010011111011111000;
	ram[841] = 58'b1000110010001111010011010111000101010111011100111011111100;
	ram[842] = 58'b1000110001111100000001001101001111010011001010010101100000;
	ram[843] = 58'b1000110001101000110000011000000000010001111101110000011101;
	ram[844] = 58'b1000110001010101100000110111010000001010101001010100000000;
	ram[845] = 58'b1000110001000010010010101010110101101111000000101000001100;
	ram[846] = 58'b1000110000101111000101110010101000010101001001111010110010;
	ram[847] = 58'b1000110000011011111010001110011111010100010110111101101001;
	ram[848] = 58'b1000110000001000101111111110010010101000000100011010110000;
	ram[849] = 58'b1000101111110101100111000001111000100011111011001110000111;
	ram[850] = 58'b1000101111100010011111011001001010001011101001110100111000;
	ram[851] = 58'b1000101111001111011001000011111101010010010100100100100101;
	ram[852] = 58'b1000101110111100010100000010001001111000000011000001101100;
	ram[853] = 58'b1000101110101001010000010011100111111110000010111010000011;
	ram[854] = 58'b1000101110010110001101111000001110100000110110110001101000;
	ram[855] = 58'b1000101110000011001100101111110101000001000111010100010000;
	ram[856] = 58'b1000101101110000001100111010010011000000100111000100101000;
	ram[857] = 58'b1000101101011101001110010111100000100101000111000000000000;
	ram[858] = 58'b1000101101001010010001000111010100001101000010101010010110;
	ram[859] = 58'b1000101100110111010101001001100110100011010001010000000000;
	ram[860] = 58'b1000101100100100011010011110001110101011010110100100000000;
	ram[861] = 58'b1000101100010001100001000101000100001100110100000011001011;
	ram[862] = 58'b1000101011111110101000111101111110110000010011111001000010;
	ram[863] = 58'b1000101011101011110010001000110101111111101000110100000100;
	ram[864] = 58'b1000101011011000111100100101100001100101101101111010000000;
	ram[865] = 58'b1000101011000110001000010011111001110001010001111111110000;
	ram[866] = 58'b1000101010110011010101010011110101001010001000100011111000;
	ram[867] = 58'b1000101010100000100011100101001100100011111010010110110100;
	ram[868] = 58'b1000101010001101110011000111110111001011010110110000011100;
	ram[869] = 58'b1000101001111011000011111011101100110001000000000111000011;
	ram[870] = 58'b1000101001101000010110000000100100100011111010110010011010;
	ram[871] = 58'b1000101001010101101001010110010111011100000011000111111001;
	ram[872] = 58'b1000101001000010111101111100111100101010101010000110000000;
	ram[873] = 58'b1000101000110000010011110100001100000100101101111001011100;
	ram[874] = 58'b1000101000011101101010111011111101100000010011001111000110;
	ram[875] = 58'b1000101000001011000011010100001000110100100101001000010101;
	ram[876] = 58'b1000100111111000011100111100100101111001110100101111010000;
	ram[877] = 58'b1000100111100101110111110101001100101001011001001011000000;
	ram[878] = 58'b1000100111010011010011111101110100111101101111010100000010;
	ram[879] = 58'b1000100111000000110001010110010110110010011001101000011001;
	ram[880] = 58'b1000100110101110001111111110101010000100000000000000000000;
	ram[881] = 58'b1000100110011011101111110110100110110000001111100000111100;
	ram[882] = 58'b1000100110001001010000111110000100110101111010010011101110;
	ram[883] = 58'b1000100101110110110011010100111100010100110111010111100101;
	ram[884] = 58'b1000100101100100010110111011000101001110000010010110110000;
	ram[885] = 58'b1000100101010001111011110000010111100011011011011010110000;
	ram[886] = 58'b1000100100111111100001110100101011011000000111000000101010;
	ram[887] = 58'b1000100100101101001001000111111000001101111100010110000100;
	ram[888] = 58'b1000100100011010110001101001110111001110101100001101001000;
	ram[889] = 58'b1000100100001000011011011010011111011100000100111001110000;
	ram[890] = 58'b1000100011110110000110011001101010000001111010010001110110;
	ram[891] = 58'b1000100011100011110010100111001110000100000110010000110100;
	ram[892] = 58'b1000100011010001100000000011000100001110010010110000010000;
	ram[893] = 58'b1000100010111111001110101101000100101010111101100100001011;
	ram[894] = 58'b1000100010101100111110100101000111100101100111011000010010;
	ram[895] = 58'b1000100010011010101111101011000101001010110011100100010000;
	ram[896] = 58'b1000100010001000100001111110110101101000001000000000000000;
	ram[897] = 58'b1000100001110110010101100000010000101010000111000000000000;
	ram[898] = 58'b1000100001100100001010001111001111000010100011010100001110;
	ram[899] = 58'b1000100001010010000000001011101001100100001101110100000000;
	ram[900] = 58'b1000100000111111110111010101010111011100101011101011111100;
	ram[901] = 58'b1000100000101101101111101100010000111110110000011100101100;
	ram[902] = 58'b1000100000011011101001010000001111100010010010100101101010;
	ram[903] = 58'b1000100000001001100100000001001010111010000001111101001001;
	ram[904] = 58'b1000011111110111011111111110111010111001110100101110111000;
	ram[905] = 58'b1000011111100101011101001001011000011010100000100100011100;
	ram[906] = 58'b1000011111010011011011100000011011110011111011100101011000;
	ram[907] = 58'b1000011111000001011011000011111100111101000001101000010100;
	ram[908] = 58'b1000011110101111011011110011110101010011100001000101000000;
	ram[909] = 58'b1000011110011101011101101111111100001110011100101111001100;
	ram[910] = 58'b1000011110001011100000111000001010101011100111010101000010;
	ram[911] = 58'b1000011101111001100101001100011000100110000010010000000000;
	ram[912] = 58'b1000011101100111101010101100011111011111010011010101110000;
	ram[913] = 58'b1000011101010101110001011000010110110010100110000011011100;
	ram[914] = 58'b1000011101000011111001001111110111100001100111101110000000;
	ram[915] = 58'b1000011100110010000010010010111001101011011100101100110100;
	ram[916] = 58'b1000011100100000001100100001010110010011101110100000101100;
	ram[917] = 58'b1000011100001110010111111011000101111101010001110101111011;
	ram[918] = 58'b1000011011111100100100100000000001001011111010000000101000;
	ram[919] = 58'b1000011011101010110010010000000000000010101011010001011001;
	ram[920] = 58'b1000011011011001000001001010111011101001000110010000101000;
	ram[921] = 58'b1000011011000111010001010000101100100101111001111111000000;
	ram[922] = 58'b1000011010110101100010100001001011100000110011011000000000;
	ram[923] = 58'b1000011010100011110100111100010000100000110100111001010000;
	ram[924] = 58'b1000011010010010001000100001110100001111101011000001000000;
	ram[925] = 58'b1000011010000000011101010001110000011011001101100100001100;
	ram[926] = 58'b1000011001101110110011001011111100001010001100100110010010;
	ram[927] = 58'b1000011001011101001010010000010001101101111110110100100100;
	ram[928] = 58'b1000011001001011100010011110101000110000111000101101100000;
	ram[929] = 58'b1000011000111001111011110110111010100010111100101000000111;
	ram[930] = 58'b1000011000101000010110011000111111110011100011101011111000;
	ram[931] = 58'b1000011000010110110010000100110000110001100011111101000101;
	ram[932] = 58'b1000011000000101001110111010000110001110010011011100000000;
	ram[933] = 58'b1000010111110011101100111000111001011101100010100110101100;
	ram[934] = 58'b1000010111100010001100000001000011010010011101010100011010;
	ram[935] = 58'b1000010111010000101100010010011100100001001011001000010001;
	ram[936] = 58'b1000010110111111001101101100111100111011111010010110000000;
	ram[937] = 58'b1000010110101101110000010000011110111100111110100110000111;
	ram[938] = 58'b1000010110011100010011111100111010011000011110011100011000;
	ram[939] = 58'b1000010110001010111000110010001000100111101011110100000000;
	ram[940] = 58'b1000010101111001011110110000000010000010000010110011010000;
	ram[941] = 58'b1000010101101000000101110110011111100001010100001011000000;
	ram[942] = 58'b1000010101010110101110000101011011000010110100111000100000;
	ram[943] = 58'b1000010101000101010111011100101011111110001011100111111001;
	ram[944] = 58'b1000010100110100000001111100001100110011110100000000000000;
	ram[945] = 58'b1000010100100010101101100011110100111101010000111100000000;
	ram[946] = 58'b1000010100010001011010010011011110111100101100100011111000;
	ram[947] = 58'b1000010100000000001000001011000010001101100101010101001101;
	ram[948] = 58'b1000010011101110110111001010011000110010100101100010101100;
	ram[949] = 58'b1000010011011101100111010001011011101100110000000000000000;
	ram[950] = 58'b1000010011001100011000100000000011011100110101001100101010;
	ram[951] = 58'b1000010010111011001010110110001001100110111001010111110001;
	ram[952] = 58'b1000010010101001111110010011100110101101100010110010001000;
	ram[953] = 58'b1000010010011000110010111000010011110101011101111011110111;
	ram[954] = 58'b1000010010000111101000100100001010100101011000011000000000;
	ram[955] = 58'b1000010001110110011111010111000100000011101101111101010100;
	ram[956] = 58'b1000010001100101010111010000111000110110101110010000000000;
	ram[957] = 58'b1000010001010100010000010001100010000110101010100100101100;
	ram[958] = 58'b1000010001000011001010011000111001011101101111101011000010;
	ram[959] = 58'b1000010000110010000101100110110111100100111011000100000000;
	ram[960] = 58'b1000010000100001000001111011010101100111000111101001000000;
	ram[961] = 58'b1000010000001111111111010110001101010001001000100100100111;
	ram[962] = 58'b1000001111111110111101110111010111001110100111010110011110;
	ram[963] = 58'b1000001111101101111101011110101101001110000101011101000000;
	ram[964] = 58'b1000001111011100111110001100000111111100111110011000011100;
	ram[965] = 58'b1000001111001011111111111111100000101010100101011001001100;
	ram[966] = 58'b1000001110111011000010111000110001001000000000001010100000;
	ram[967] = 58'b1000001110101010000110110111110010000101010100001110000100;
	ram[968] = 58'b1000001110011001001011111100011101010101010011110111111000;
	ram[969] = 58'b1000001110001000010010000110101011001000111110000100100111;
	ram[970] = 58'b1000001101110111011001010110010110010110100001010100010110;
	ram[971] = 58'b1000001101100110100001101011010110101111110110001111110100;
	ram[972] = 58'b1000001101010101101011000101100110101011111110010011010000;
	ram[973] = 58'b1000001101000100110101100100111111000000001111101010001100;
	ram[974] = 58'b1000001100110100000001001001011001000011101101001111001000;
	ram[975] = 58'b1000001100100011001101110010101110101111000001110110011001;
	ram[976] = 58'b1000001100010010011011100000111000111010001001101100000000;
	ram[977] = 58'b1000001100000001101010010011110001011111011001100101011100;
	ram[978] = 58'b1000001011110000111010001011010000110111101110011110111110;
	ram[979] = 58'b1000001011100000001011000111010001011111110110110001001101;
	ram[980] = 58'b1000001011001111011101000111101100010011001010110101001100;
	ram[981] = 58'b1000001010111110110000001100011011001111010010011101001100;
	ram[982] = 58'b1000001010101110000100010101010110110000101001011010100000;
	ram[983] = 58'b1000001010011101011001100010011001010111001011111111010001;
	ram[984] = 58'b1000001010001100101111110011011100000001101100001010100000;
	ram[985] = 58'b1000001001111100000111001000011000110001000010110011011100;
	ram[986] = 58'b1000001001101011011111100001001000000101001000000001100110;
	ram[987] = 58'b1000001001011010111000111101100100100001000100001101010101;
	ram[988] = 58'b1000001001001010010011011101100111000111000000101110000100;
	ram[989] = 58'b1000001000111001101111000001001001111011000101001110101100;
	ram[990] = 58'b1000001000101001001011101000000101100000100100100001001000;
	ram[991] = 58'b1000001000011000101001010010010100011101110000011101101001;
	ram[992] = 58'b1000001000001000000111111111101111111000001000000000000000;
	ram[993] = 58'b1000000111110111100111110000010001010110100000110101011111;
	ram[994] = 58'b1000000111100111001000100011110010100000100100011100111000;
	ram[995] = 58'b1000000111010110101010011010001101011111001100110100000000;
	ram[996] = 58'b1000000111000110001101010011011011011011001100000001110000;
	ram[997] = 58'b1000000110110101110001001111010101011110001100011010111011;
	ram[998] = 58'b1000000110100101010110001101110110010011111011011100001010;
	ram[999] = 58'b1000000110010100111100001110110111101000000001000000000000;
	ram[1000] = 58'b1000000110000100100011010010010010000110001001110001100000;
	ram[1001] = 58'b1000000101110100001011010111111111111100000000000000000000;
	ram[1002] = 58'b1000000101100011110100011111111011010111111101000010110110;
	ram[1003] = 58'b1000000101010011011110101001111101101000100000001110010100;
	ram[1004] = 58'b1000000101000011001001110101111111111101000000000000000000;
	ram[1005] = 58'b1000000100110010110110000011111101000110011111011000001011;
	ram[1006] = 58'b1000000100100010100011010011101110010101111000011000001000;
	ram[1007] = 58'b1000000100010010010001100101001101011101001011011011101001;
	ram[1008] = 58'b1000000100000010000000111000010100101111011010010110010000;
	ram[1009] = 58'b1000000011110001110001001100111100111111101010010111000000;
	ram[1010] = 58'b1000000011100001100010100011000000100010100001110111001110;
	ram[1011] = 58'b1000000011010001010100111010011001101101010101011011000101;
	ram[1012] = 58'b1000000011000001001000010011000001110101110000010110101100;
	ram[1013] = 58'b1000000010110000111100101100110010010010010100010110101100;
	ram[1014] = 58'b1000000010100000110010000111100101111010110010110111101000;
	ram[1015] = 58'b1000000010010000101000100011010110000111001110110101100100;
	ram[1016] = 58'b1000000010000000011111111111111100010000100000011100001000;
	ram[1017] = 58'b1000000001110000011000011101010011010000100110110110001111;
	ram[1018] = 58'b1000000001100000010001111011010100100001111010111100110110;
	ram[1019] = 58'b1000000001010000001100011001111001111111101110100011010101;
	ram[1020] = 58'b1000000001000000000111111000111101100110000100000111000100;
	ram[1021] = 58'b1000000000110000000100011000011001010001101110100111111011;
	ram[1022] = 58'b1000000000100000000001111000000111000000010001100000110010;
	ram[1023] = 58'b1000000000010000000000011000000000110000000000100000000001;
end
endmodule

module finv_load_grad_table (
    input wire [9:0] addr,
    output wire [34:0] grd,
    input wire clk,
	input wire rstn);

(* RAM_STYLE="BLOCK" *) reg [34:0] ram [1023:0];
//always @(posedge clk)
//    grd <= ram[addr];
assign grd = ram[addr];
initial begin
	ram[0] = 35'b11111111110000000001001111111110000;
	ram[1] = 35'b11111111010000000111001111100010000;
	ram[2] = 35'b11111110110000010011001101111110001;
	ram[3] = 35'b11111110010000100101000010100100010;
	ram[4] = 35'b11111101110000111100111100100001111;
	ram[5] = 35'b11111101010001011010100011001101110;
	ram[6] = 35'b11111100110001111110001101110001111;
	ram[7] = 35'b11111100010010100111100011101000100;
	ram[8] = 35'b11111011110011010110110011111100101;
	ram[9] = 35'b11111011010100001011111101111111001;
	ram[10] = 35'b11111010110101000110110001001011001;
	ram[11] = 35'b11111010010110000111010100101111000;
	ram[12] = 35'b11111001110111001101101111110110111;
	ram[13] = 35'b11111001011000011001110010000001001;
	ram[14] = 35'b11111000111001101011100010011011000;
	ram[15] = 35'b11111000011011000011000000010111000;
	ram[16] = 35'b11110111111100100000000011010000001;
	ram[17] = 35'b11110111011110000010101010011010111;
	ram[18] = 35'b11110110111111101011000100111001011;
	ram[19] = 35'b11110110100001011000111010011010000;
	ram[20] = 35'b11110110000011001100011001111110110;
	ram[21] = 35'b11110101100101000101011011000101100;
	ram[22] = 35'b11110101000111000011111101000011000;
	ram[23] = 35'b11110100101001000111111111001100000;
	ram[24] = 35'b11110100001011010001011001000001101;
	ram[25] = 35'b11110011101101100000011001100001010;
	ram[26] = 35'b11110011001111110100110000011000100;
	ram[27] = 35'b11110010110010001110100100110000101;
	ram[28] = 35'b11110010010100101101110101111110111;
	ram[29] = 35'b11110001110111010010011011100111000;
	ram[30] = 35'b11110001011001111100010100111111111;
	ram[31] = 35'b11110000111100101011101001010001000;
	ram[32] = 35'b11110000011111100000010000000000000;
	ram[33] = 35'b11110000000010011010001000100011101;
	ram[34] = 35'b11101111100101011001010010010011011;
	ram[35] = 35'b11101111001000011101101100100110011;
	ram[36] = 35'b11101110101011100111010110110011111;
	ram[37] = 35'b11101110001110110110010000010011011;
	ram[38] = 35'b11101101110010001010010000101110111;
	ram[39] = 35'b11101101010101100011011111001100011;
	ram[40] = 35'b11101100111001000001111011000011011;
	ram[41] = 35'b11101100011100100101011011111111101;
	ram[42] = 35'b11101100000000001110001001000101111;
	ram[43] = 35'b11101011100011111011111010000010111;
	ram[44] = 35'b11101011000111101110101110001111111;
	ram[45] = 35'b11101010101011100110100101000110010;
	ram[46] = 35'b11101010001111100011100101101001011;
	ram[47] = 35'b11101001110011100101011111111110101;
	ram[48] = 35'b11101001010111101100100010110010110;
	ram[49] = 35'b11101000111011111000011110001101011;
	ram[50] = 35'b11101000100000001001011001010001011;
	ram[51] = 35'b11101000000100011111001011110001001;
	ram[52] = 35'b11100111101000111010000100010110000;
	ram[53] = 35'b11100111001101011001110011001011011;
	ram[54] = 35'b11100110110001111110010111101100110;
	ram[55] = 35'b11100110010110100111111000111011001;
	ram[56] = 35'b11100101111011010110001110101011101;
	ram[57] = 35'b11100101100000001001011000011001101;
	ram[58] = 35'b11100101000101000001010101100000111;
	ram[59] = 35'b11100100101001111110001101000001001;
	ram[60] = 35'b11100100001110111111101111001101110;
	ram[61] = 35'b11100011110100000110001010101001111;
	ram[62] = 35'b11100011011001010001001111101011010;
	ram[63] = 35'b11100010111110100001000101010001001;
	ram[64] = 35'b11100010100011110101101010110111101;
	ram[65] = 35'b11100010001001001110111000011001110;
	ram[66] = 35'b11100001101110101100111100010110010;
	ram[67] = 35'b11100001010100001111011111100111011;
	ram[68] = 35'b11100000111001110110110000101011110;
	ram[69] = 35'b11100000011111100010100111100000011;
	ram[70] = 35'b11100000000101010011001011000001111;
	ram[71] = 35'b11011111101011001000010011001110011;
	ram[72] = 35'b11011111010001000001111111100011110;
	ram[73] = 35'b11011110110111000000001111011111110;
	ram[74] = 35'b11011110011101000011000010100000101;
	ram[75] = 35'b11011110000011001010010000100111100;
	ram[76] = 35'b11011101101001010110001000001100101;
	ram[77] = 35'b11011101001111100110100001010001000;
	ram[78] = 35'b11011100110101111011010011110111010;
	ram[79] = 35'b11011100011100010100100110111010010;
	ram[80] = 35'b11011100000010110010010010011101100;
	ram[81] = 35'b11011011101001010100011101011011010;
	ram[82] = 35'b11011011001111111011000111010001110;
	ram[83] = 35'b11011010110110100110000000101101000;
	ram[84] = 35'b11011010011101010101011000000000000;
	ram[85] = 35'b11011010000100001001001100101001011;
	ram[86] = 35'b11011001101011000001001111010111110;
	ram[87] = 35'b11011001010001111101101110011011111;
	ram[88] = 35'b11011000111000111110011010100110001;
	ram[89] = 35'b11011000100000000011100010000101100;
	ram[90] = 35'b11011000000111001100110101101100011;
	ram[91] = 35'b11010111101110011010011100010010001;
	ram[92] = 35'b11010111010101101100010101010111001;
	ram[93] = 35'b11010110111101000010100000011011111;
	ram[94] = 35'b11010110100100011100110101101100010;
	ram[95] = 35'b11010110001011111011011011111110001;
	ram[96] = 35'b11010101110011011110001011011110010;
	ram[97] = 35'b11010101011011000101001011000010010;
	ram[98] = 35'b11010101000010110000010010110111011;
	ram[99] = 35'b11010100101010011111100010100000000;
	ram[100] = 35'b11010100010010010011000000110000010;
	ram[101] = 35'b11010011111010001010100101110111001;
	ram[102] = 35'b11010011100010000110010001010111000;
	ram[103] = 35'b11010011001010000110000010110010000;
	ram[104] = 35'b11010010110010001001110010011001101;
	ram[105] = 35'b11010010011010010001101110010010001;
	ram[106] = 35'b11010010000010011101101110101100101;
	ram[107] = 35'b11010001101010101101101011111100011;
	ram[108] = 35'b11010001010011000001101100110100000;
	ram[109] = 35'b11010000111011011001110000110110000;
	ram[110] = 35'b11010000100011110101110111100101000;
	ram[111] = 35'b11010000001100010101110010001000001;
	ram[112] = 35'b11001111110100111001110101101100101;
	ram[113] = 35'b11001111011101100001110011011010000;
	ram[114] = 35'b11001111000110001101101010110100011;
	ram[115] = 35'b11001110101110111101011011011111111;
	ram[116] = 35'b11001110010111110001001100001100010;
	ram[117] = 35'b11001110000000101000110101010001001;
	ram[118] = 35'b11001101101001100100010110010010111;
	ram[119] = 35'b11001101010010100011100111101011000;
	ram[120] = 35'b11001100111011100110110111010011011;
	ram[121] = 35'b11001100100100101101111101100101011;
	ram[122] = 35'b11001100001101111000111010000101101;
	ram[123] = 35'b11001011110111000111100101001111011;
	ram[124] = 35'b11001011100000011010001100111001100;
	ram[125] = 35'b11001011001001110000100010010111001;
	ram[126] = 35'b11001010110011001010100101001110000;
	ram[127] = 35'b11001010011100101000011100001011011;
	ram[128] = 35'b11001010000110001010000110110011110;
	ram[129] = 35'b11001001101111101111011101100101101;
	ram[130] = 35'b11001001011001011000100000000110110;
	ram[131] = 35'b11001001000011000101010101000010111;
	ram[132] = 35'b11001000101100110101110100111001101;
	ram[133] = 35'b11001000010110101001111111010001001;
	ram[134] = 35'b11001000000000100001111010110100000;
	ram[135] = 35'b11000111101010011101011000111111000;
	ram[136] = 35'b11000111010100011100100111100001001;
	ram[137] = 35'b11000110111110011111010111111000100;
	ram[138] = 35'b11000110101000100101110111110011000;
	ram[139] = 35'b11000110010010101111111000110000010;
	ram[140] = 35'b11000101111100111101100001011010001;
	ram[141] = 35'b11000101100111001110110001010111010;
	ram[142] = 35'b11000101010001100011101000001110001;
	ram[143] = 35'b11000100111011111011111110100100000;
	ram[144] = 35'b11000100100110010111111011000001100;
	ram[145] = 35'b11000100010000110111010110001100111;
	ram[146] = 35'b11000011111011011010010110101110000;
	ram[147] = 35'b11000011100110000000110101001011111;
	ram[148] = 35'b11000011010000101010111000001101101;
	ram[149] = 35'b11000010111011011000011000011011011;
	ram[150] = 35'b11000010100110001001010101011101000;
	ram[151] = 35'b11000010010000111101110101111000101;
	ram[152] = 35'b11000001111011110101101011011001111;
	ram[153] = 35'b11000001100110110001000011100100101;
	ram[154] = 35'b11000001010001101111110111000010111;
	ram[155] = 35'b11000000111100110010000101011101000;
	ram[156] = 35'b11000000100111110111100111011110111;
	ram[157] = 35'b11000000010011000000101010101001100;
	ram[158] = 35'b10111111111110001101000000101101011;
	ram[159] = 35'b10111111101001011100110000001111000;
	ram[160] = 35'b10111111010100101111111000110110110;
	ram[161] = 35'b10111111000000000110011010001101000;
	ram[162] = 35'b10111110101011100000001101000000011;
	ram[163] = 35'b10111110010110111101010111110100000;
	ram[164] = 35'b10111110000010011101110011010111011;
	ram[165] = 35'b10111101101110000001100110001100111;
	ram[166] = 35'b10111101011001101000101001000100111;
	ram[167] = 35'b10111101000101010011000010100001000;
	ram[168] = 35'b10111100110001000000100100011010111;
	ram[169] = 35'b10111100011100110001100011000011001;
	ram[170] = 35'b10111100001000100101101001011100111;
	ram[171] = 35'b10111011110100011100111110001001100;
	ram[172] = 35'b10111011100000010111100111101001011;
	ram[173] = 35'b10111011001100010101011110101111011;
	ram[174] = 35'b10111010111000010110011100010000010;
	ram[175] = 35'b10111010100100011010101101100001011;
	ram[176] = 35'b10111010010000100010000100100010001;
	ram[177] = 35'b10111001111100101100101110100110101;
	ram[178] = 35'b10111001101000111010011101110000000;
	ram[179] = 35'b10111001010101001011011000011101001;
	ram[180] = 35'b10111001000001011111011110011000010;
	ram[181] = 35'b10111000101101110110101000011000111;
	ram[182] = 35'b10111000011010010000111100111100111;
	ram[183] = 35'b10111000000110101110010100111100011;
	ram[184] = 35'b10110111110011001110110110110100111;
	ram[185] = 35'b10110111011111110010100010010000101;
	ram[186] = 35'b10110111001100011001010000001001001;
	ram[187] = 35'b10110110111001000011000000001001111;
	ram[188] = 35'b10110110100101101111111000101111000;
	ram[189] = 35'b10110110010010011111110010110011000;
	ram[190] = 35'b10110101111111010010101110000001100;
	ram[191] = 35'b10110101101100001000101010000110010;
	ram[192] = 35'b10110101011001000001100110101101000;
	ram[193] = 35'b10110101000101111101101010010000010;
	ram[194] = 35'b10110100110010111100100110111110001;
	ram[195] = 35'b10110100011111111110101001111111011;
	ram[196] = 35'b10110100001101000011100101100011110;
	ram[197] = 35'b10110011111010001011100110110010110;
	ram[198] = 35'b10110011100111010110011111111101010;
	ram[199] = 35'b10110011010100100100010111011101001;
	ram[200] = 35'b10110011000001110101001100111110010;
	ram[201] = 35'b10110010101111001000111001100000110;
	ram[202] = 35'b10110010011100011111101010001000111;
	ram[203] = 35'b10110010001001111001001010100000011;
	ram[204] = 35'b10110001110111010101101110010101101;
	ram[205] = 35'b10110001100100110101000111111111000;
	ram[206] = 35'b10110001010010010111010111001001110;
	ram[207] = 35'b10110000111111111100100010001100111;
	ram[208] = 35'b10110000101101100100100010001011011;
	ram[209] = 35'b10110000011011001111011101011011100;
	ram[210] = 35'b10110000001000111101001101000001000;
	ram[211] = 35'b10101111110110101101110000101001001;
	ram[212] = 35'b10101111100100100001001000000001100;
	ram[213] = 35'b10101111010010010111011001011111001;
	ram[214] = 35'b10101111000000010000011110000111010;
	ram[215] = 35'b10101110101110001100001111000000011;
	ram[216] = 35'b10101110011100001010111001000110011;
	ram[217] = 35'b10101110001010001100010101011111100;
	ram[218] = 35'b10101101111000010000100011111001010;
	ram[219] = 35'b10101101100110010111011101011011111;
	ram[220] = 35'b10101101010100100001001111000000100;
	ram[221] = 35'b10101101000010101101101011001010000;
	ram[222] = 35'b10101100110000111100111110110000010;
	ram[223] = 35'b10101100011111001110110101110011001;
	ram[224] = 35'b10101100001101100011100011101110100;
	ram[225] = 35'b10101011111011111010111011000111110;
	ram[226] = 35'b10101011101010010101000010010001001;
	ram[227] = 35'b10101011011000110001111000111000011;
	ram[228] = 35'b10101011000111010001011000001001000;
	ram[229] = 35'b10101010110101110011011111110001111;
	ram[230] = 35'b10101010100100011000010110000011111;
	ram[231] = 35'b10101010010010111111110100001011010;
	ram[232] = 35'b10101010000001101010000000011000101;
	ram[233] = 35'b10101001110000010110110011111000110;
	ram[234] = 35'b10101001011111000110001110011011000;
	ram[235] = 35'b10101001001101111000010110001110101;
	ram[236] = 35'b10101000111100101100111110000001111;
	ram[237] = 35'b10101000101011100100010010100100001;
	ram[238] = 35'b10101000011010011110001101000100010;
	ram[239] = 35'b10101000001001011010101101010001100;
	ram[240] = 35'b10100111111000011001110010111011010;
	ram[241] = 35'b10100111100111011011100100001110111;
	ram[242] = 35'b10100111010110011111110011111110110;
	ram[243] = 35'b10100111000101100110101000011000111;
	ram[244] = 35'b10100110110100101111111010101111011;
	ram[245] = 35'b10100110100011111011110111101100011;
	ram[246] = 35'b10100110010011001010010010000101001;
	ram[247] = 35'b10100110000010011011010110100010100;
	ram[248] = 35'b10100101110001101110110111111011010;
	ram[249] = 35'b10100101100001000100110101111111101;
	ram[250] = 35'b10100101010000011101010110111011100;
	ram[251] = 35'b10100100111111111000011010011110011;
	ram[252] = 35'b10100100101111010110000000010111110;
	ram[253] = 35'b10100100011110110110000001111101000;
	ram[254] = 35'b10100100001110011000011110111110100;
	ram[255] = 35'b10100011111101111101011101100110101;
	ram[256] = 35'b10100011101101100100110111001011101;
	ram[257] = 35'b10100011011101001110110001110111011;
	ram[258] = 35'b10100011001100111011000111000000101;
	ram[259] = 35'b10100010111100101001110110011000001;
	ram[260] = 35'b10100010101100011010111111101110100;
	ram[261] = 35'b10100010011100001110101001001100100;
	ram[262] = 35'b10100010001100000100101100001010010;
	ram[263] = 35'b10100001111011111101001000011000101;
	ram[264] = 35'b10100001101011110111111101101000011;
	ram[265] = 35'b10100001011011110101001011101010011;
	ram[266] = 35'b10100001001011110100110010001111011;
	ram[267] = 35'b10100000111011110110110001001000011;
	ram[268] = 35'b10100000101011111011001000000110010;
	ram[269] = 35'b10100000011100000001110110111001111;
	ram[270] = 35'b10100000001100001010111101010100010;
	ram[271] = 35'b10011111111100010110011011000110011;
	ram[272] = 35'b10011111101100100100010000000001001;
	ram[273] = 35'b10011111011100110100010101100001100;
	ram[274] = 35'b10011111001101000110110001101101011;
	ram[275] = 35'b10011110111101011011100100010101100;
	ram[276] = 35'b10011110101101110010100110111000001;
	ram[277] = 35'b10011110011110001011111111011010000;
	ram[278] = 35'b10011110001110100111101101101100010;
	ram[279] = 35'b10011101111111000101101011001101110;
	ram[280] = 35'b10011101101111100101111110000010101;
	ram[281] = 35'b10011101100000001000011111101010100;
	ram[282] = 35'b10011101010000101101001111110111011;
	ram[283] = 35'b10011101000001010100010100101100100;
	ram[284] = 35'b10011100110001111101101101111011010;
	ram[285] = 35'b10011100100010101001001110110011111;
	ram[286] = 35'b10011100010011010111000011101001111;
	ram[287] = 35'b10011100000100000111001100001110101;
	ram[288] = 35'b10011011110100111001011011110100011;
	ram[289] = 35'b10011011100101101101111110101100111;
	ram[290] = 35'b10011011010110100100101110011010100;
	ram[291] = 35'b10011011000111011101101010101111101;
	ram[292] = 35'b10011010111000011000110011011110100;
	ram[293] = 35'b10011010101001010110001000011001110;
	ram[294] = 35'b10011010011010010101101001010011101;
	ram[295] = 35'b10011010001011010111010101111110101;
	ram[296] = 35'b10011001111100011011001110001101000;
	ram[297] = 35'b10011001101101100001010001110001011;
	ram[298] = 35'b10011001011110101001100000011110010;
	ram[299] = 35'b10011001001111110011111010000110000;
	ram[300] = 35'b10011001000001000000011110011011010;
	ram[301] = 35'b10011000110010001111000111000101000;
	ram[302] = 35'b10011000100011011111111010000001111;
	ram[303] = 35'b10011000010100110010110111000100011;
	ram[304] = 35'b10011000000110000111110111110100110;
	ram[305] = 35'b10010111110111011111001000011011000;
	ram[306] = 35'b10010111101000111000010110001010101;
	ram[307] = 35'b10010111011010010011110011010101101;
	ram[308] = 35'b10010111001011110001010011011010101;
	ram[309] = 35'b10010110111101010000110110001101011;
	ram[310] = 35'b10010110101110110010100001101010001;
	ram[311] = 35'b10010110100000010110010101100100000;
	ram[312] = 35'b10010110010001111100001011100101001;
	ram[313] = 35'b10010110000011100100000011100001010;
	ram[314] = 35'b10010101110101001101111101001100001;
	ram[315] = 35'b10010101100110111001111110100000111;
	ram[316] = 35'b10010101011000101000000111010010010;
	ram[317] = 35'b10010101001010011000001011000101100;
	ram[318] = 35'b10010100111100001010010101111100011;
	ram[319] = 35'b10010100101101111110100001100011011;
	ram[320] = 35'b10010100011111110100101101101110100;
	ram[321] = 35'b10010100010001101100111010010001100;
	ram[322] = 35'b10010100000011100111000111000000001;
	ram[323] = 35'b10010011110101100011011001110011010;
	ram[324] = 35'b10010011100111100001100110010100100;
	ram[325] = 35'b10010011011001100001111000100001011;
	ram[326] = 35'b10010011001011100100000100000100110;
	ram[327] = 35'b10010010111101101000010100111011000;
	ram[328] = 35'b10010010101111101110011110110000001;
	ram[329] = 35'b10010010100001110110100111011100010;
	ram[330] = 35'b10010010010100000000101110110011010;
	ram[331] = 35'b10010010000110001100110100101001001;
	ram[332] = 35'b10010001111000011010111000110010000;
	ram[333] = 35'b10010001101010101010110100111111100;
	ram[334] = 35'b10010001011100111100101111001000101;
	ram[335] = 35'b10010001001111010000100111000001011;
	ram[336] = 35'b10010001000001100110011100011101111;
	ram[337] = 35'b10010000110011111110001001010001000;
	ram[338] = 35'b10010000100110010111110011010000101;
	ram[339] = 35'b10010000011000110011010100010000011;
	ram[340] = 35'b10010000001011010000110010000101011;
	ram[341] = 35'b10001111111101110000001100100011111;
	ram[342] = 35'b10001111110000010001011101100000011;
	ram[343] = 35'b10001111100010110100100100101111111;
	ram[344] = 35'b10001111010101011001101000000110100;
	ram[345] = 35'b10001111001000000000100111011000110;
	ram[346] = 35'b10001110111010101001010110011101011;
	ram[347] = 35'b10001110101101010100000001000111010;
	ram[348] = 35'b10001110100000000000100111001010011;
	ram[349] = 35'b10001110010010101110111100011111110;
	ram[350] = 35'b10001110000101011111001100111000001;
	ram[351] = 35'b10001101111000010001010010001010111;
	ram[352] = 35'b10001101101011000101010010001001111;
	ram[353] = 35'b10001101011101111011000000110000100;
	ram[354] = 35'b10001101010000110010101001101101001;
	ram[355] = 35'b10001101000011101100000000111100011;
	ram[356] = 35'b10001100110110100111010010001011110;
	ram[357] = 35'b10001100101001100100010111010100001;
	ram[358] = 35'b10001100011100100011010000001010111;
	ram[359] = 35'b10001100001111100011111100100101001;
	ram[360] = 35'b10001100000010100110011100011000100;
	ram[361] = 35'b10001011110101101010101111011010000;
	ram[362] = 35'b10001011101000110000110101011111001;
	ram[363] = 35'b10001011011011111000101000100011011;
	ram[364] = 35'b10001011001111000010010100010000001;
	ram[365] = 35'b10001011000010001101101100100111001;
	ram[366] = 35'b10001010110101011010110111010111111;
	ram[367] = 35'b10001010101000101001110100010111110;
	ram[368] = 35'b10001010011011111010100011011100001;
	ram[369] = 35'b10001010001111001101000100011010011;
	ram[370] = 35'b10001010000010100001010001010000010;
	ram[371] = 35'b10001001110101110111001001110011110;
	ram[372] = 35'b10001001101001001110111001101010001;
	ram[373] = 35'b10001001011100101000010100111001110;
	ram[374] = 35'b10001001010000000011100001010000000;
	ram[375] = 35'b10001001000011100000011000101011101;
	ram[376] = 35'b10001000110110111111000000111001010;
	ram[377] = 35'b10001000101010011111010011111000101;
	ram[378] = 35'b10001000011110000001010111010101110;
	ram[379] = 35'b10001000010001100101000101010000110;
	ram[380] = 35'b10001000000101001010011101100000000;
	ram[381] = 35'b10000111111000110001101011100100000;
	ram[382] = 35'b10000111101100011010011101110011011;
	ram[383] = 35'b10000111100000000100111111101110010;
	ram[384] = 35'b10000111010011110001001011010110000;
	ram[385] = 35'b10000111000111011111000000100001011;
	ram[386] = 35'b10000110111011001110100100111010010;
	ram[387] = 35'b10000110101110111111110010100011010;
	ram[388] = 35'b10000110100010110010101001010010100;
	ram[389] = 35'b10000110010110100111001000111110111;
	ram[390] = 35'b10000110001010011101010111010001011;
	ram[391] = 35'b10000101111110010101001000011011001;
	ram[392] = 35'b10000101110010001110100111110111101;
	ram[393] = 35'b10000101100110001001101111101010111;
	ram[394] = 35'b10000101011010000110011111101011011;
	ram[395] = 35'b10000101001110000100110001111110100;
	ram[396] = 35'b10000101000010000100110001111101111;
	ram[397] = 35'b10000100110110000110011001101110011;
	ram[398] = 35'b10000100101010001001101001000110111;
	ram[399] = 35'b10000100011110001110011111111101110;
	ram[400] = 35'b10000100010010010100111110001001111;
	ram[401] = 35'b10000100000110011100111101110010001;
	ram[402] = 35'b10000011111010100110101010001101000;
	ram[403] = 35'b10000011101110110001110111110010000;
	ram[404] = 35'b10000011100010111110101100000111100;
	ram[405] = 35'b10000011010111001101000111000100010;
	ram[406] = 35'b10000011001011011101001000011111010;
	ram[407] = 35'b10000010111111101110101010100000110;
	ram[408] = 35'b10000010110100000001110010101110011;
	ram[409] = 35'b10000010101000010110100000111110111;
	ram[410] = 35'b10000010011100101100110101001001001;
	ram[411] = 35'b10000010010001000100101001010110110;
	ram[412] = 35'b10000010000101011101111101011111011;
	ram[413] = 35'b10000001111001111000111100110011111;
	ram[414] = 35'b10000001101110010101011011110001101;
	ram[415] = 35'b10000001100010110011011010010000000;
	ram[416] = 35'b10000001010111010010111101110010111;
	ram[417] = 35'b10000001001011110100000110010001000;
	ram[418] = 35'b10000001000000010110101000001010100;
	ram[419] = 35'b10000000110100111010110100011001010;
	ram[420] = 35'b10000000101001100000011111011101100;
	ram[421] = 35'b10000000011110000111101001001111010;
	ram[422] = 35'b10000000010010110000010001100101111;
	ram[423] = 35'b10000000000111011010011110000011100;
	ram[424] = 35'b01111111111100000110001000110101001;
	ram[425] = 35'b01111111110000110011010111011100001;
	ram[426] = 35'b01111111100101100010000100000110001;
	ram[427] = 35'b01111111011010010010001110101010111;
	ram[428] = 35'b01111111001111000011110111000010010;
	ram[429] = 35'b01111111000011110111000010101100100;
	ram[430] = 35'b01111110111000101011101011111000100;
	ram[431] = 35'b01111110101101100001101100110101110;
	ram[432] = 35'b01111110100010011001010110010100110;
	ram[433] = 35'b01111110010111010010010111010100101;
	ram[434] = 35'b01111110001100001100110101010101100;
	ram[435] = 35'b01111110000001001000110000001111001;
	ram[436] = 35'b01111101110110000110001101100000100;
	ram[437] = 35'b01111101101011000101000001110011010;
	ram[438] = 35'b01111101100000000101010010100110100;
	ram[439] = 35'b01111101010101000111000101011000011;
	ram[440] = 35'b01111101001010001010001110110100000;
	ram[441] = 35'b01111100111111001110111001111101101;
	ram[442] = 35'b01111100110100010100111011100001100;
	ram[443] = 35'b01111100101001011100011000111101100;
	ram[444] = 35'b01111100011110100101010010001001100;
	ram[445] = 35'b01111100010011101111100110111101101;
	ram[446] = 35'b01111100001000111011010001101101001;
	ram[447] = 35'b01111011111110001000011101011001101;
	ram[448] = 35'b01111011110011010110111110110010000;
	ram[449] = 35'b01111011101000100110111011010010111;
	ram[450] = 35'b01111011011101111000010010110100011;
	ram[451] = 35'b01111011010011001010111111101011001;
	ram[452] = 35'b01111011001000011111001100110110001;
	ram[453] = 35'b01111010111101110100101001100100000;
	ram[454] = 35'b01111010110011001011100110010110011;
	ram[455] = 35'b01111010101000100011110111111111101;
	ram[456] = 35'b01111010011101111101100011111010111;
	ram[457] = 35'b01111010010011011000100100011110001;
	ram[458] = 35'b01111010001000110100111111000100000;
	ram[459] = 35'b01111001111110010010101110000011010;
	ram[460] = 35'b01111001110011110001110110110101110;
	ram[461] = 35'b01111001101001010010011001010011110;
	ram[462] = 35'b01111001011110110100001111110100101;
	ram[463] = 35'b01111001010100010111011010010001011;
	ram[464] = 35'b01111001001001111011111110000011000;
	ram[465] = 35'b01111000111111100001110101100001111;
	ram[466] = 35'b01111000110101001001000110000110011;
	ram[467] = 35'b01111000101010110001101010001001011;
	ram[468] = 35'b01111000100000011011100001100011110;
	ram[469] = 35'b01111000010110000110110001101101100;
	ram[470] = 35'b01111000001011110011010101000000000;
	ram[471] = 35'b01111000000001100001010000110010111;
	ram[472] = 35'b01110111110111010000011010000001101;
	ram[473] = 35'b01110111101101000000111011100010010;
	ram[474] = 35'b01110111100010110010101111101111000;
	ram[475] = 35'b01110111011000100101110110100000111;
	ram[476] = 35'b01110111001110011010010101001110011;
	ram[477] = 35'b01110111000100010000000110010010101;
	ram[478] = 35'b01110110111010000111000100001001110;
	ram[479] = 35'b01110110101111111111011001100110110;
	ram[480] = 35'b01110110100101111001000001000101100;
	ram[481] = 35'b01110110011011110011111111111011100;
	ram[482] = 35'b01110110010001110000001011001000111;
	ram[483] = 35'b01110110000111101101101000000011010;
	ram[484] = 35'b01110101111101101100010110100011101;
	ram[485] = 35'b01110101110011101100011011111110100;
	ram[486] = 35'b01110101101001101101101101010110000;
	ram[487] = 35'b01110101011111110000001111111110111;
	ram[488] = 35'b01110101010101110100000011110010010;
	ram[489] = 35'b01110101001011111001001110000011100;
	ram[490] = 35'b01110101000001111111100011110110111;
	ram[491] = 35'b01110100111000000111001010100000000;
	ram[492] = 35'b01110100101110001111111100011110011;
	ram[493] = 35'b01110100100100011010000100011110111;
	ram[494] = 35'b01110100011010100101011101000000110;
	ram[495] = 35'b01110100010000110010000000100100000;
	ram[496] = 35'b01110100000110111111110100011011011;
	ram[497] = 35'b01110011111101001110111000100000000;
	ram[498] = 35'b01110011110011011111001100101011001;
	ram[499] = 35'b01110011101001110000101011011101111;
	ram[500] = 35'b01110011100000000011011010001010000;
	ram[501] = 35'b01110011010110010111011000101000110;
	ram[502] = 35'b01110011001100101100100001011011111;
	ram[503] = 35'b01110011000011000010111001110100100;
	ram[504] = 35'b01110010111001011010100001101100000;
	ram[505] = 35'b01110010101111110011011000111011101;
	ram[506] = 35'b01110010100110001101011010000101111;
	ram[507] = 35'b01110010011100101000100101000101000;
	ram[508] = 35'b01110010010011000100111111001000111;
	ram[509] = 35'b01110010001001100010101000001010110;
	ram[510] = 35'b01110010000000000001011010101110100;
	ram[511] = 35'b01110001110110100001011100000011011;
	ram[512] = 35'b01110001101101000010100110101101100;
	ram[513] = 35'b01110001100011100100111111111100000;
	ram[514] = 35'b01110001011010001000100010010011010;
	ram[515] = 35'b01110001010000101101010011000001111;
	ram[516] = 35'b01110001000111010011001100101101000;
	ram[517] = 35'b01110000111101111010001111001110100;
	ram[518] = 35'b01110000110100100010011111110100100;
	ram[519] = 35'b01110000101011001011111001000100101;
	ram[520] = 35'b01110000100001110110011010111000111;
	ram[521] = 35'b01110000011000100010001010011110100;
	ram[522] = 35'b01110000001111001111000010011100001;
	ram[523] = 35'b01110000000101111101000111111110011;
	ram[524] = 35'b01101111111100101100010000011001101;
	ram[525] = 35'b01101111110011011100100110001101011;
	ram[526] = 35'b01101111101010001110000100000000111;
	ram[527] = 35'b01101111100001000000101111000000010;
	ram[528] = 35'b01101111010111110100011100100001011;
	ram[529] = 35'b01101111001110101001010111000010010;
	ram[530] = 35'b01101111000101011111011001001010110;
	ram[531] = 35'b01101110111100010110100010110101011;
	ram[532] = 35'b01101110110011001110110011111100000;
	ram[533] = 35'b01101110101010001000010001101001100;
	ram[534] = 35'b01101110100001000010110001010110101;
	ram[535] = 35'b01101110010111111110011101011110100;
	ram[536] = 35'b01101110001110111011001011011010101;
	ram[537] = 35'b01101110000101111001000101100101101;
	ram[538] = 35'b01101101111100111000000001011001101;
	ram[539] = 35'b01101101110011111000001001010000011;
	ram[540] = 35'b01101101101010111001010111110100010;
	ram[541] = 35'b01101101100001111011100111110000011;
	ram[542] = 35'b01101101011000111111000011011101011;
	ram[543] = 35'b01101101010000000011100000010111100;
	ram[544] = 35'b01101101000111001001001000110110011;
	ram[545] = 35'b01101100111110001111110010010111011;
	ram[546] = 35'b01101100110101010111100010000011011;
	ram[547] = 35'b01101100101100100000010111110100100;
	ram[548] = 35'b01101100100011101010010011100101001;
	ram[549] = 35'b01101100011010110101010101001111011;
	ram[550] = 35'b01101100010010000001010111100000110;
	ram[551] = 35'b01101100001001001110100100101101100;
	ram[552] = 35'b01101100000000011100110010010110010;
	ram[553] = 35'b01101011110111101100000101100010011;
	ram[554] = 35'b01101011101110111100011110001100000;
	ram[555] = 35'b01101011100110001101110111000001101;
	ram[556] = 35'b01101011011101100000010101001010000;
	ram[557] = 35'b01101011010100110011111000011111010;
	ram[558] = 35'b01101011001100001000100000111011111;
	ram[559] = 35'b01101011000011011110001001001111001;
	ram[560] = 35'b01101010111010110100110110011110110;
	ram[561] = 35'b01101010110010001100100011011010100;
	ram[562] = 35'b01101010101001100101010101000111111;
	ram[563] = 35'b01101010100000111111001011100001001;
	ram[564] = 35'b01101010011000011010000001010110110;
	ram[565] = 35'b01101010001111110101111011101101011;
	ram[566] = 35'b01101010000111010010111010011111101;
	ram[567] = 35'b01101001111110110000110011010101000;
	ram[568] = 35'b01101001110110001111110101100100101;
	ram[569] = 35'b01101001101101101111110110110110100;
	ram[570] = 35'b01101001100101010000110111000101100;
	ram[571] = 35'b01101001011100110010111011010101011;
	ram[572] = 35'b01101001010100010110000011100000100;
	ram[573] = 35'b01101001001011111010001010011001010;
	ram[574] = 35'b01101001000011011111001111111010100;
	ram[575] = 35'b01101000111011000101011001000111010;
	ram[576] = 35'b01101000110010101100100000110010010;
	ram[577] = 35'b01101000101010010100100110110110110;
	ram[578] = 35'b01101000100001111101110000010110111;
	ram[579] = 35'b01101000011001100111111000000110010;
	ram[580] = 35'b01101000010001010011000011000110101;
	ram[581] = 35'b01101000001000111111001100001100001;
	ram[582] = 35'b01101000000000101100010011010001101;
	ram[583] = 35'b01100111111000011010011000010010011;
	ram[584] = 35'b01100111110000001001100000001111100;
	ram[585] = 35'b01100111100111111001100101111101110;
	ram[586] = 35'b01100111011111101010101001011000001;
	ram[587] = 35'b01100111010111011100101111011111010;
	ram[588] = 35'b01100111001111001111101110000011011;
	ram[589] = 35'b01100111000111000011101111001010010;
	ram[590] = 35'b01100110111110111000101101101001011;
	ram[591] = 35'b01100110110110101110101110100000110;
	ram[592] = 35'b01100110101110100101100111100010010;
	ram[593] = 35'b01100110100110011101011101101101101;
	ram[594] = 35'b01100110011110010110010110000010001;
	ram[595] = 35'b01100110010110010000001011010110101;
	ram[596] = 35'b01100110001110001010111000100010110;
	ram[597] = 35'b01100110000110000110100111101000111;
	ram[598] = 35'b01100101111110000011010011100000101;
	ram[599] = 35'b01100101110110000000111100000101010;
	ram[600] = 35'b01100101101101111111100001010001110;
	ram[601] = 35'b01100101100101111111000011000001101;
	ram[602] = 35'b01100101011101111111100001001111111;
	ram[603] = 35'b01100101010110000000111011110111111;
	ram[604] = 35'b01100101001110000011010010110100111;
	ram[605] = 35'b01100101000110000110100110000010000;
	ram[606] = 35'b01100100111110001010110101011010101;
	ram[607] = 35'b01100100110110010000000000111010001;
	ram[608] = 35'b01100100101110010110000011011010011;
	ram[609] = 35'b01100100100110011101000110111001010;
	ram[610] = 35'b01100100011110100101000110010000110;
	ram[611] = 35'b01100100010110101101111100011011100;
	ram[612] = 35'b01100100001110110111101110010101110;
	ram[613] = 35'b01100100000111000010011011111010111;
	ram[614] = 35'b01100011111111001110000101000110001;
	ram[615] = 35'b01100011110111011010101001110010111;
	ram[616] = 35'b01100011101111101000000100111100110;
	ram[617] = 35'b01100011100111110110011011011111010;
	ram[618] = 35'b01100011100000000101101101010101011;
	ram[619] = 35'b01100011011000010101111010011010110;
	ram[620] = 35'b01100011010000100111000010101010101;
	ram[621] = 35'b01100011001000111001000001000001101;
	ram[622] = 35'b01100011000001001011111010011010010;
	ram[623] = 35'b01100010111001011111101110101111110;
	ram[624] = 35'b01100010110001110100011000111111100;
	ram[625] = 35'b01100010101010001001111110000011010;
	ram[626] = 35'b01100010100010100000011101110110011;
	ram[627] = 35'b01100010011010110111110011010110111;
	ram[628] = 35'b01100010010011010000000011011110000;
	ram[629] = 35'b01100010001011101001001001001001111;
	ram[630] = 35'b01100010000100000011001110010000100;
	ram[631] = 35'b01100001111100011110000011110110011;
	ram[632] = 35'b01100001110100111001111000101101101;
	ram[633] = 35'b01100001101101010110100010111000101;
	ram[634] = 35'b01100001100101110100000010010011001;
	ram[635] = 35'b01100001011110010010011011110101001;
	ram[636] = 35'b01100001010110110001101010011110100;
	ram[637] = 35'b01100001001111010001110011000110101;
	ram[638] = 35'b01100001000111110010110101101000111;
	ram[639] = 35'b01100001000000010100101101000101110;
	ram[640] = 35'b01100000111000110111011001011001001;
	ram[641] = 35'b01100000110001011010111111011001110;
	ram[642] = 35'b01100000101001111111011010001000101;
	ram[643] = 35'b01100000100010100100101110011100001;
	ram[644] = 35'b01100000011011001010110111010101100;
	ram[645] = 35'b01100000010011110001111001101010111;
	ram[646] = 35'b01100000001100011001110000011101110;
	ram[647] = 35'b01100000000101000010011011101010011;
	ram[648] = 35'b01011111111101101100000000000110001;
	ram[649] = 35'b01011111110110010110011000110011010;
	ram[650] = 35'b01011111101111000001100101101101111;
	ram[651] = 35'b01011111100111101101100110110010001;
	ram[652] = 35'b01011111100000011010100000110100101;
	ram[653] = 35'b01011111011001001000010011110000111;
	ram[654] = 35'b01011111010001110110110101110001111;
	ram[655] = 35'b01011111001010100110010000100100101;
	ram[656] = 35'b01011111000011010110011111001100100;
	ram[657] = 35'b01011110111100000111100001100101101;
	ram[658] = 35'b01011110110100111001011100100011111;
	ram[659] = 35'b01011110101101101100000110010011110;
	ram[660] = 35'b01011110100110011111101000100000101;
	ram[661] = 35'b01011110011111010011111110001110110;
	ram[662] = 35'b01011110011000001001001100010001011;
	ram[663] = 35'b01011110010000111111001000110110100;
	ram[664] = 35'b01011110001001110101111101100111111;
	ram[665] = 35'b01011110000010101101100000110100100;
	ram[666] = 35'b01011101111011100101111100000101010;
	ram[667] = 35'b01011101110100011111001010011111111;
	ram[668] = 35'b01011101101101011001001100000000011;
	ram[669] = 35'b01011101100110010100000000100011001;
	ram[670] = 35'b01011101011111001111101100111001100;
	ram[671] = 35'b01011101011000001100000111010100101;
	ram[672] = 35'b01011101010001001001010100100110100;
	ram[673] = 35'b01011101001010000111011001011111111;
	ram[674] = 35'b01011101000011000110001100010011010;
	ram[675] = 35'b01011100111100000101110001110001110;
	ram[676] = 35'b01011100110101000110001110101011111;
	ram[677] = 35'b01011100101110000111011001010101001;
	ram[678] = 35'b01011100100111001001011011010001111;
	ram[679] = 35'b01011100100000001100001010110110100;
	ram[680] = 35'b01011100011001001111101100110011001;
	ram[681] = 35'b01011100010010010100000001000100010;
	ram[682] = 35'b01011100001011011001001100011001000;
	ram[683] = 35'b01011100000100011111000101000111001;
	ram[684] = 35'b01011011111101100101101111111110001;
	ram[685] = 35'b01011011110110101101001000000111110;
	ram[686] = 35'b01011011101111110101010111000101101;
	ram[687] = 35'b01011011101000111110011000000001001;
	ram[688] = 35'b01011011100010001000000110000100100;
	ram[689] = 35'b01011011011011010010101010110000010;
	ram[690] = 35'b01011011010100011101111100011100101;
	ram[691] = 35'b01011011001101101001111111111000000;
	ram[692] = 35'b01011011000110110110110000001101001;
	ram[693] = 35'b01011011000000000100010110111011011;
	ram[694] = 35'b01011010111001010010101010011100100;
	ram[695] = 35'b01011010110010100001101111011101111;
	ram[696] = 35'b01011010101011110001100101111100000;
	ram[697] = 35'b01011010100101000010001101110011000;
	ram[698] = 35'b01011010011110010011100010001111000;
	ram[699] = 35'b01011010010111100101100111111100110;
	ram[700] = 35'b01011010010000111000011110111000110;
	ram[701] = 35'b01011010001010001100000010001111011;
	ram[702] = 35'b01011010000011100000011011011100110;
	ram[703] = 35'b01011001111100110101011100001110010;
	ram[704] = 35'b01011001110110001011010010101111010;
	ram[705] = 35'b01011001101111100001110101011101000;
	ram[706] = 35'b01011001101000111001001001000011101;
	ram[707] = 35'b01011001100010010001001000110000011;
	ram[708] = 35'b01011001011011101001111001001110111;
	ram[709] = 35'b01011001010101000011011010011011011;
	ram[710] = 35'b01011001001110011101100111100100000;
	ram[711] = 35'b01011001000111111000100101010011110;
	ram[712] = 35'b01011001000001010100001110111000111;
	ram[713] = 35'b01011000111010110000101000111110010;
	ram[714] = 35'b01011000110100001101110011100000000;
	ram[715] = 35'b01011000101101101011101001101101001;
	ram[716] = 35'b01011000100111001010001011100010101;
	ram[717] = 35'b01011000100000101001100010010111011;
	ram[718] = 35'b01011000011010001001100000000000100;
	ram[719] = 35'b01011000010011101010001101110101000;
	ram[720] = 35'b01011000001101001011101011110001010;
	ram[721] = 35'b01011000000110101101110101000101001;
	ram[722] = 35'b01011000000000010000101001101101101;
	ram[723] = 35'b01010111111001110100001110010011110;
	ram[724] = 35'b01010111110011011000100010110011101;
	ram[725] = 35'b01010111101100111101100010011110010;
	ram[726] = 35'b01010111100110100011001101010000011;
	ram[727] = 35'b01010111100000001001100011000111000;
	ram[728] = 35'b01010111011001110000101101010101011;
	ram[729] = 35'b01010111010011011000011101110110011;
	ram[730] = 35'b01010111001101000000111101111101000;
	ram[731] = 35'b01010111000110101010001000111011010;
	ram[732] = 35'b01010111000000010011111110101101111;
	ram[733] = 35'b01010110111001111110100011111100010;
	ram[734] = 35'b01010110110011101001110011111000100;
	ram[735] = 35'b01010110101101010101110011001001110;
	ram[736] = 35'b01010110100111000010011101000010011;
	ram[737] = 35'b01010110100000101111110001011111101;
	ram[738] = 35'b01010110011010011101110000011110011;
	ram[739] = 35'b01010110010100001100011110100100101;
	ram[740] = 35'b01010110001101111011110111000110001;
	ram[741] = 35'b01010110000111101011111001111111100;
	ram[742] = 35'b01010110000001011100101011110110101;
	ram[743] = 35'b01010101111011001110000011010110110;
	ram[744] = 35'b01010101110101000000001001101110010;
	ram[745] = 35'b01010101101110110010111010010001011;
	ram[746] = 35'b01010101101000100110010100111101000;
	ram[747] = 35'b01010101100010011010011110010110000;
	ram[748] = 35'b01010101011100001111010001110001011;
	ram[749] = 35'b01010101010110000100101010100100010;
	ram[750] = 35'b01010101001111111010110001111011001;
	ram[751] = 35'b01010101001001110001100111110010011;
	ram[752] = 35'b01010101000011101001000010111000100;
	ram[753] = 35'b01010100111101100001000111110001110;
	ram[754] = 35'b01010100110111011001111011000010000;
	ram[755] = 35'b01010100110001010011010111111111001;
	ram[756] = 35'b01010100101011001101011001111111110;
	ram[757] = 35'b01010100100101001000001010001101111;
	ram[758] = 35'b01010100011111000011100100000000000;
	ram[759] = 35'b01010100011000111111100111010011001;
	ram[760] = 35'b01010100010010111100010100000100010;
	ram[761] = 35'b01010100001100111001101010010000011;
	ram[762] = 35'b01010100000110110111101001110100101;
	ram[763] = 35'b01010100000000110110010010101110000;
	ram[764] = 35'b01010011111010110101101001011110110;
	ram[765] = 35'b01010011110100110101100100111001011;
	ram[766] = 35'b01010011101110110110001001100000010;
	ram[767] = 35'b01010011101000110111010111010000100;
	ram[768] = 35'b01010011100010111001001110000111001;
	ram[769] = 35'b01010011011100111011101110000001010;
	ram[770] = 35'b01010011010110111110110110111011110;
	ram[771] = 35'b01010011010001000010101000110100000;
	ram[772] = 35'b01010011001011000111000011100110110;
	ram[773] = 35'b01010011000101001100000111010001011;
	ram[774] = 35'b01010010111111010001110011110000101;
	ram[775] = 35'b01010010111001011000000100011110101;
	ram[776] = 35'b01010010110011011111000010011110111;
	ram[777] = 35'b01010010101101100110100100101000011;
	ram[778] = 35'b01010010100111101110110011111110001;
	ram[779] = 35'b01010010100001110111100111010111011;
	ram[780] = 35'b01010010011100000001000011010100010;
	ram[781] = 35'b01010010010110001011000111110010000;
	ram[782] = 35'b01010010010000010101110100101101100;
	ram[783] = 35'b01010010001010100001000101100010000;
	ram[784] = 35'b01010010000100101101000011010000110;
	ram[785] = 35'b01010001111110111001100100110011000;
	ram[786] = 35'b01010001111001000110101110100111111;
	ram[787] = 35'b01010001110011010100100000101100100;
	ram[788] = 35'b01010001101101100010110110011100110;
	ram[789] = 35'b01010001100111110001111000111000011;
	ram[790] = 35'b01010001100010000001011110111010001;
	ram[791] = 35'b01010001011100010001101101000000101;
	ram[792] = 35'b01010001010110100010011110101000001;
	ram[793] = 35'b01010001010000110011111000001110110;
	ram[794] = 35'b01010001001011000101111001110001110;
	ram[795] = 35'b01010001000101011000100011001110001;
	ram[796] = 35'b01010000111111101011110100100001010;
	ram[797] = 35'b01010000111001111111101001001000001;
	ram[798] = 35'b01010000110100010100000101100000011;
	ram[799] = 35'b01010000101110101001000101000111011;
	ram[800] = 35'b01010000101000111110101100011010011;
	ram[801] = 35'b01010000100011010100111011010110010;
	ram[802] = 35'b01010000011101101011110001111000011;
	ram[803] = 35'b01010000011000000011001011011111000;
	ram[804] = 35'b01010000010010011011001100100110100;
	ram[805] = 35'b01010000001100110011110000101101011;
	ram[806] = 35'b01010000000111001100111100001111110;
	ram[807] = 35'b01010000000001100110101111001010111;
	ram[808] = 35'b01001111111100000001000100111101110;
	ram[809] = 35'b01001111110110011100000010000100000;
	ram[810] = 35'b01001111110000110111100001111101001;
	ram[811] = 35'b01001111101011010011101001000100010;
	ram[812] = 35'b01001111100101110000010010111001001;
	ram[813] = 35'b01001111100000001101100011110110111;
	ram[814] = 35'b01001111011010101011011011111010101;
	ram[815] = 35'b01001111010101001001110110100100100;
	ram[816] = 35'b01001111001111101000111000001111000;
	ram[817] = 35'b01001111001010001000011100011010111;
	ram[818] = 35'b01001111000100101000100011000101101;
	ram[819] = 35'b01001110111111001001010000101001011;
	ram[820] = 35'b01001110111001101010100101000011010;
	ram[821] = 35'b01001110110100001100011011110100100;
	ram[822] = 35'b01001110101110101110111001010110110;
	ram[823] = 35'b01001110101001010001111001001011011;
	ram[824] = 35'b01001110100011110101011011010000010;
	ram[825] = 35'b01001110011110011001100011111110010;
	ram[826] = 35'b01001110011000111110001110110111100;
	ram[827] = 35'b01001110010011100011100000010100110;
	ram[828] = 35'b01001110001110001001010011111000011;
	ram[829] = 35'b01001110001000101111101101111010111;
	ram[830] = 35'b01001110000011010110101001111110110;
	ram[831] = 35'b01001101111101111110001000000001110;
	ram[832] = 35'b01001101111000100110001100011100000;
	ram[833] = 35'b01001101110011001110110010110000100;
	ram[834] = 35'b01001101101101110111111010111101000;
	ram[835] = 35'b01001101101000100001101001011001001;
	ram[836] = 35'b01001101100011001011111001101000011;
	ram[837] = 35'b01001101011101110110110000000010001;
	ram[838] = 35'b01001101011000100010001000001010001;
	ram[839] = 35'b01001101010011001110000001111110001;
	ram[840] = 35'b01001101001101111010011101011011110;
	ram[841] = 35'b01001101001000100111011110111010000;
	ram[842] = 35'b01001101000011010101000001111101001;
	ram[843] = 35'b01001100111110000011000110100010111;
	ram[844] = 35'b01001100111000110001110001000001110;
	ram[845] = 35'b01001100110011100000111100111110010;
	ram[846] = 35'b01001100101110010000101010010110100;
	ram[847] = 35'b01001100101001000000111001001000000;
	ram[848] = 35'b01001100100011110001101101101000101;
	ram[849] = 35'b01001100011110100010111111000101111;
	ram[850] = 35'b01001100011001010100111010100101010;
	ram[851] = 35'b01001100010100000111010010111100110;
	ram[852] = 35'b01001100001110111010001100100010001;
	ram[853] = 35'b01001100001001101101101011101010010;
	ram[854] = 35'b01001100000100100001101011111011100;
	ram[855] = 35'b01001011111111010110001101010011101;
	ram[856] = 35'b01001011111010001011001111110000010;
	ram[857] = 35'b01001011110101000000110111100110000;
	ram[858] = 35'b01001011101111110110111100000101001;
	ram[859] = 35'b01001011101010101101100101111000100;
	ram[860] = 35'b01001011100101100100110000100111010;
	ram[861] = 35'b01001011100000011100011100001111010;
	ram[862] = 35'b01001011011011010100101000101110010;
	ram[863] = 35'b01001011010110001101010110000010000;
	ram[864] = 35'b01001011010001000110100100001000011;
	ram[865] = 35'b01001011001100000000010111010100101;
	ram[866] = 35'b01001011000110111010100110111001011;
	ram[867] = 35'b01001011000001110101011011011111010;
	ram[868] = 35'b01001010111100110000110000101110101;
	ram[869] = 35'b01001010110111101100100110100101010;
	ram[870] = 35'b01001010110010101000111000101100010;
	ram[871] = 35'b01001010101101100101101111101011000;
	ram[872] = 35'b01001010101000100011000111001010011;
	ram[873] = 35'b01001010100011100000111111001000011;
	ram[874] = 35'b01001010011110011111010111100010101;
	ram[875] = 35'b01001010011001011110010000010111000;
	ram[876] = 35'b01001010010100011101101001100011011;
	ram[877] = 35'b01001010001111011101100011000101100;
	ram[878] = 35'b01001010001010011101111100111011010;
	ram[879] = 35'b01001010000101011110110111000010100;
	ram[880] = 35'b01001010000000100000010001011001000;
	ram[881] = 35'b01001001111011100010001011111100100;
	ram[882] = 35'b01001001110110100100100110101011000;
	ram[883] = 35'b01001001110001100111100001100010001;
	ram[884] = 35'b01001001101100101010111100100000000;
	ram[885] = 35'b01001001100111101110110111100010010;
	ram[886] = 35'b01001001100010110011010010100110110;
	ram[887] = 35'b01001001011101111000001001011001001;
	ram[888] = 35'b01001001011000111101100100011011111;
	ram[889] = 35'b01001001010100000011011011001000100;
	ram[890] = 35'b01001001001111001001110110000000111;
	ram[891] = 35'b01001001001010010000101100011111001;
	ram[892] = 35'b01001001000101011000000010110011000;
	ram[893] = 35'b01001001000000011111111000111010011;
	ram[894] = 35'b01001000111011101000001110110011001;
	ram[895] = 35'b01001000110110110001000100011011001;
	ram[896] = 35'b01001000110001111010011001110000010;
	ram[897] = 35'b01001000101101000100001010011111100;
	ram[898] = 35'b01001000101000001110011010110111111;
	ram[899] = 35'b01001000100011011001001111000111111;
	ram[900] = 35'b01001000011110100100011110101011111;
	ram[901] = 35'b01001000011001110000001001100010100;
	ram[902] = 35'b01001000010100111100011000001010001;
	ram[903] = 35'b01001000010000001001000110010000010;
	ram[904] = 35'b01001000001011010110001111100010111;
	ram[905] = 35'b01001000000110100011111000010000001;
	ram[906] = 35'b01001000000001110010000000010101110;
	ram[907] = 35'b01000111111101000000100011100010010;
	ram[908] = 35'b01000111111000001111101010010010101;
	ram[909] = 35'b01000111110011011111001100000101111;
	ram[910] = 35'b01000111101110101111001101001001100;
	ram[911] = 35'b01000111101001111111101001001100011;
	ram[912] = 35'b01000111100101010000101000101010011;
	ram[913] = 35'b01000111100000100010000011000011110;
	ram[914] = 35'b01000111011011110011111100100101010;
	ram[915] = 35'b01000111010111000110010000111110100;
	ram[916] = 35'b01000111010010011001000100011100001;
	ram[917] = 35'b01000111001101101100010110111011111;
	ram[918] = 35'b01000111001001000000001000011011110;
	ram[919] = 35'b01000111000100010100010100101011110;
	ram[920] = 35'b01000110111111101000111111111000001;
	ram[921] = 35'b01000110111010111110001001111110100;
	ram[922] = 35'b01000110110110010011110010111100111;
	ram[923] = 35'b01000110110001101001110110100100001;
	ram[924] = 35'b01000110101101000000010100110010011;
	ram[925] = 35'b01000110101000010111010110000000000;
	ram[926] = 35'b01000110100011101110101101100100000;
	ram[927] = 35'b01000110011111000110101000000011001;
	ram[928] = 35'b01000110011010011110111101000001111;
	ram[929] = 35'b01000110010101110111110000101011001;
	ram[930] = 35'b01000110010001010001000010111100101;
	ram[931] = 35'b01000110001100101010101111101000010;
	ram[932] = 35'b01000110001000000100110110101100011;
	ram[933] = 35'b01000110000011011111011100010011010;
	ram[934] = 35'b01000101111110111010100000011010110;
	ram[935] = 35'b01000101111010010110000011000000110;
	ram[936] = 35'b01000101110101110001111011101100100;
	ram[937] = 35'b01000101110001001110010110111110100;
	ram[938] = 35'b01000101101100101011001100011110001;
	ram[939] = 35'b01000101101000001000100000010100110;
	ram[940] = 35'b01000101100011100110001110010101010;
	ram[941] = 35'b01000101011111000100010110011110010;
	ram[942] = 35'b01000101011010100011000001000011010;
	ram[943] = 35'b01000101010110000010000001100010011;
	ram[944] = 35'b01000101010001100001100100011001011;
	ram[945] = 35'b01000101001101000001011101000111010;
	ram[946] = 35'b01000101001000100001111000001000111;
	ram[947] = 35'b01000101000100000010101000111110010;
	ram[948] = 35'b01000100111111100011110111111001101;
	ram[949] = 35'b01000100111011000101100100111001000;
	ram[950] = 35'b01000100110110100111101011110000110;
	ram[951] = 35'b01000100110010001010010000101000110;
	ram[952] = 35'b01000100101101101101001111010101101;
	ram[953] = 35'b01000100101001010000100111110101111;
	ram[954] = 35'b01000100100100110100011110010000111;
	ram[955] = 35'b01000100100000011000110010100100100;
	ram[956] = 35'b01000100011011111101100000100110001;
	ram[957] = 35'b01000100010111100010101000010100001;
	ram[958] = 35'b01000100010011001000001101110101010;
	ram[959] = 35'b01000100001110101110001100111111011;
	ram[960] = 35'b01000100001010010100100101110000110;
	ram[961] = 35'b01000100000101111011011100001111111;
	ram[962] = 35'b01000100000001100010101100010010111;
	ram[963] = 35'b01000011111101001010011001111111111;
	ram[964] = 35'b01000011111000110010100001001101010;
	ram[965] = 35'b01000011110100011011000001111001011;
	ram[966] = 35'b01000011110000000100000000001010001;
	ram[967] = 35'b01000011101011101101010111110110001;
	ram[968] = 35'b01000011100111010111001101000011001;
	ram[969] = 35'b01000011100011000001010111100001000;
	ram[970] = 35'b01000011011110101100000011100011001;
	ram[971] = 35'b01000011011010010111000100110011000;
	ram[972] = 35'b01000011010110000010100011011100110;
	ram[973] = 35'b01000011010001101110011011010111101;
	ram[974] = 35'b01000011001101011010101100100010011;
	ram[975] = 35'b01000011001001000111011011000001100;
	ram[976] = 35'b01000011000100110100100010101100111;
	ram[977] = 35'b01000011000000100010000111101001000;
	ram[978] = 35'b01000010111100010000000001101000001;
	ram[979] = 35'b01000010110111111110011000110100101;
	ram[980] = 35'b01000010110011101101001001000110111;
	ram[981] = 35'b01000010101111011100010110100010111;
	ram[982] = 35'b01000010101011001011111000111011111;
	ram[983] = 35'b01000010100110111011111000011011000;
	ram[984] = 35'b01000010100010101100010000111001100;
	ram[985] = 35'b01000010011110011101000110011010101;
	ram[986] = 35'b01000010011010001110010000110010111;
	ram[987] = 35'b01000010010101111111111000001010010;
	ram[988] = 35'b01000010010001110001111000011010100;
	ram[989] = 35'b01000010001101100100010101100110011;
	ram[990] = 35'b01000010001001010111000111100011010;
	ram[991] = 35'b01000010000101001010010110011000100;
	ram[992] = 35'b01000010000000111101111110000000000;
	ram[993] = 35'b01000001111100110001111110011000010;
	ram[994] = 35'b01000001111000100110010111011111101;
	ram[995] = 35'b01000001110100011011001101011000011;
	ram[996] = 35'b01000001110000010000011011111101000;
	ram[997] = 35'b01000001101100000101111111001000100;
	ram[998] = 35'b01000001100111111011111111000000011;
	ram[999] = 35'b01000001100011110010011011100010100;
	ram[1000] = 35'b01000001011111101001001100100111001;
	ram[1001] = 35'b01000001011011100000010110010000000;
	ram[1002] = 35'b01000001010111010111111100011110001;
	ram[1003] = 35'b01000001010011001111111011001101001;
	ram[1004] = 35'b01000001001111001000001110011001000;
	ram[1005] = 35'b01000001001011000000111110000101001;
	ram[1006] = 35'b01000001000110111010000110001101101;
	ram[1007] = 35'b01000001000010110011100110110000111;
	ram[1008] = 35'b01000000111110101101100011101111010;
	ram[1009] = 35'b01000000111010100111110101000011001;
	ram[1010] = 35'b01000000110110100010011110101101010;
	ram[1011] = 35'b01000000110010011101100100101101101;
	ram[1012] = 35'b01000000101110011001000011000000111;
	ram[1013] = 35'b01000000101010010100110101100100001;
	ram[1014] = 35'b01000000100110010001000100011000101;
	ram[1015] = 35'b01000000100010001101101011011011011;
	ram[1016] = 35'b01000000011110001010100110101010001;
	ram[1017] = 35'b01000000011010000111111110000101001;
	ram[1018] = 35'b01000000010110000101101101101001111;
	ram[1019] = 35'b01000000010010000011110101010111000;
	ram[1020] = 35'b01000000001110000010010101001010111;
	ram[1021] = 35'b01000000001010000001001101000100000;
	ram[1022] = 35'b01000000000110000000011101000000111;
	ram[1023] = 35'b01000000000010000000000101000000000;
end
endmodule
`default_nettype wire