`timescale 1ns / 100ps
`default_nettype none

module test_itof
    #(parameter NSTAGE = 2,
      parameter REPEATNUM = 50,
      parameter RANDSEED = 2) ();

wire [31:0] x1,y;
shortreal    fx1, fy, absfy;
logic [31:0] absx, fybit, absfybit;

logic clk, rstn;
int i, diff;
logic [31:0] r, x1d;

logic [31:0] x1_reg[NSTAGE:0];
logic val[NSTAGE:0];

assign x1 = x1_reg[0];

itof u1(x1,y,clk,rstn);

initial begin
	// $dumpfile("test_itof.vcd");
	// $dumpvars(0);

    $display("start of checking module itof");
    $display("difference message format");
    $display("x1 = [input 1(bit)], [exponent 1(decimal)]");
    $display("x2 = [input 2(bit)], [exponent 2(decimal)]");
    $display("ref. : result(float) sign(bit),exponent(decimal),mantissa(bit)");
    $display("itof : result(float) sign(bit),exponent(decimal),mantissa(bit)");
    
    #1;			//t = 1ns
    rstn = 0;
    clk = 1;
    val = {default: 1'b0};
    x1_reg[0] = 0;
    i=0;

    #1;			//t = 2ns
    clk = 0;
    #1;			//t = 3ns
    clk = 1;
    rstn = 1;

    repeat(RANDSEED) begin
        i = $urandom();
    end

    repeat(REPEATNUM) begin
        r = $urandom();
        x1d = $urandom();
        x1_reg[0] <= (r[0]) ? x1d : {x1d[31], 21'b0, x1d[9:0]};
        val[0] <= 1;

        #1;
		clk = 0;
		#1;
		clk = 1;
        /*
        repeat(NSTAGE) begin
            #1;
		    clk = 0;
		    #1;
		    clk = 1;
            val[0] <= 0;
        end
        */
    end
    repeat(NSTAGE+1) begin
        #1;
	    clk = 0;
	    #1;
	    clk = 1;
    end
    $display("end of checking module itof");
    $finish;
end

always @(posedge clk) begin
	x1_reg[NSTAGE:1] <= x1_reg[NSTAGE-1:0];
	val[NSTAGE:1] <= val[NSTAGE-1:0];
end
   
always @(posedge clk) begin
	if (val[NSTAGE]) begin      //ここ、ステージ分けがちゃんとしていれば別に必要ないです。
		
        absx = (x1_reg[NSTAGE][31] == 1) ? (~x1_reg[NSTAGE]) + 1 : x1_reg[NSTAGE];
        absfy = $itor(absx);
        absfybit = $shortrealtobits(absfy);
        fybit = {x1_reg[NSTAGE][31], absfybit[30:0]};
        fy = $bitstoshortreal(fybit);

        diff = (fybit >= y) ? fybit - y : y - fybit;
        $display("diff = %d", diff);
        //if(diff >= 1) begin
   	        $display("x = %b, %d",
	        x1_reg[NSTAGE], $signed(x1_reg[NSTAGE]));
   	        $display("%.15f %b,%3d,%b", fy,
	        fybit[31], fybit[30:23], fybit[22:0]);
   	        $display("%.15f %b,%3d,%b\n", $bitstoshortreal(y),
	        y[31], y[30:23], y[22:0]);
        //end
    end
    //$display("val = %b, %b, %b", val[0], val[1], val[2]);
    //$display("%e %b,%3d,%b %b\n", $bitstoshortreal(y),y[31], y[30:23], y[22:0], ovf);
end
endmodule

`default_nettype wire
