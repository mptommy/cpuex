`default_nettype none
module floor #(parameter NSTAGE = 2)(
    input wire [31:0] x,
    output wire [31:0] y,
    input wire clk,
    input wire rstn);

// stage = 0 (x)

// stage = 1 (xr[0] -> mni, restbit, xep)

reg [31:0] xr[1:0];

wire [7:0] e = xr[0][30:23];
wire [22:0] m = xr[0][22:0];

wire [23:0] mni =   (e <= 8'b01111111) ? 24'b0 :
                    (e == 8'b10000000) ? {1'b0, m[22], 22'b0} :
                    (e == 8'b10000001) ? {1'b0, m[22:21], 21'b0} :
                    (e == 8'b10000010) ? {1'b0, m[22:20], 20'b0} :
                    (e == 8'b10000011) ? {1'b0, m[22:19], 19'b0} :
                    (e == 8'b10000100) ? {1'b0, m[22:18], 18'b0} :
                    (e == 8'b10000101) ? {1'b0, m[22:17], 17'b0} :
                    (e == 8'b10000110) ? {1'b0, m[22:16], 16'b0} :
                    (e == 8'b10000111) ? {1'b0, m[22:15], 15'b0} :
                    (e == 8'b10001000) ? {1'b0, m[22:14], 14'b0} :
                    (e == 8'b10001001) ? {1'b0, m[22:13], 13'b0} :
                    (e == 8'b10001010) ? {1'b0, m[22:12], 12'b0} :
                    (e == 8'b10001011) ? {1'b0, m[22:11], 11'b0} :
                    (e == 8'b10001100) ? {1'b0, m[22:10], 10'b0} :
                    (e == 8'b10001101) ? {1'b0, m[22:9], 9'b0} :
                    (e == 8'b10001110) ? {1'b0, m[22:8], 8'b0} :
                    (e == 8'b10001111) ? {1'b0, m[22:7], 7'b0} :
                    (e == 8'b10010000) ? {1'b0, m[22:6], 6'b0} :
                    (e == 8'b10010001) ? {1'b0, m[22:5], 5'b0} :
                    (e == 8'b10010010) ? {1'b0, m[22:4], 4'b0} :
                    (e == 8'b10010011) ? {1'b0, m[22:3], 3'b0} :
                    (e == 8'b10010100) ? {1'b0, m[22:2], 2'b0} :
                    (e == 8'b10010101) ? {1'b0, m[22:1], 1'b0} : {1'b0, m};

wire [23:0] restbit =   (e <= 8'b01111111) ? {|(m[22:0]), 23'b0} :
                        (e == 8'b10000000) ? {1'b0, |(m[21:0]), 22'b0} :
                        (e == 8'b10000001) ? {2'b0, |(m[20:0]), 21'b0} :
                        (e == 8'b10000010) ? {3'b0, |(m[19:0]), 20'b0} :
                        (e == 8'b10000011) ? {4'b0, |(m[18:0]), 19'b0} :
                        (e == 8'b10000100) ? {5'b0, |(m[17:0]), 18'b0} :
                        (e == 8'b10000101) ? {6'b0, |(m[16:0]), 17'b0} :
                        (e == 8'b10000110) ? {7'b0, |(m[15:0]), 16'b0} :
                        (e == 8'b10000111) ? {8'b0, |(m[14:0]), 15'b0} :
                        (e == 8'b10001000) ? {9'b0, |(m[13:0]), 14'b0} :
                        (e == 8'b10001001) ? {10'b0, |(m[12:0]), 13'b0} :
                        (e == 8'b10001010) ? {11'b0, |(m[11:0]), 12'b0} :
                        (e == 8'b10001011) ? {12'b0, |(m[10:0]), 11'b0} :
                        (e == 8'b10001100) ? {13'b0, |(m[9:0]), 10'b0} :
                        (e == 8'b10001101) ? {14'b0, |(m[8:0]), 9'b0} :
                        (e == 8'b10001110) ? {15'b0, |(m[7:0]), 8'b0} :
                        (e == 8'b10001111) ? {16'b0, |(m[6:0]), 7'b0} :
                        (e == 8'b10010000) ? {17'b0, |(m[5:0]), 6'b0} :
                        (e == 8'b10010001) ? {18'b0, |(m[4:0]), 5'b0} :
                        (e == 8'b10010010) ? {19'b0, |(m[3:0]), 4'b0} :
                        (e == 8'b10010011) ? {20'b0, |(m[2:0]), 3'b0} :
                        (e == 8'b10010100) ? {21'b0, |(m[1:0]), 2'b0} :
                        (e == 8'b10010101) ? {22'b0, m[0], 1'b0} : 24'b0;

wire [7:0] xep = (e < 8'b01111111) ? 8'b0 : e;

// stage = 2 (mnir, restbitr, xepr -> y)

reg [31:0] mnir;
reg [23:0] restbitr;
reg [7:0] xepr;

wire ys = xr[1][31];

wire [23:0] mp = (ys) ? mnir + restbitr : mnir;

wire [8:0] ep = (xepr == 8'b0) ? ((mp[23]) ? 9'b001111111 : 9'b000000000) : xepr + mp[23];

wire [7:0] ye = ep[7:0];
wire [22:0] ym = (mp[23]) ? {1'b0, mp[22:1]} : mp[22:0];

always @(posedge clk) begin
    if(~rstn) begin
        xr[0] <= 'b0;
        mnir <= 'b0;
        restbitr <= 'b0;
        xepr <= 'b0;
    end else begin
        xr[0] <= x;
        mnir <= mni;
        restbitr <= restbit;
        xepr <= xep;
    end
end

always @(posedge clk) begin
    xr[1] <= xr[0];
end

assign y = {ys, ye, ym};

endmodule
`default_nettype wire